library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity applemouse_rom is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(10 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of applemouse_rom is
	type rom is array(0 to  2047) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"2C",X"58",X"FF",X"70",X"1B",X"38",X"90",X"18",X"B8",X"50",X"15",X"01",X"20",X"F4",X"F4",X"F4",
		X"F4",X"00",X"B3",X"C4",X"9B",X"A4",X"C0",X"8A",X"DD",X"BC",X"48",X"F0",X"53",X"E1",X"E6",X"EC",
		X"08",X"78",X"8D",X"F8",X"07",X"48",X"98",X"48",X"8A",X"48",X"20",X"58",X"FF",X"BA",X"BD",X"00",
		X"01",X"AA",X"08",X"0A",X"0A",X"0A",X"0A",X"28",X"A8",X"AD",X"F8",X"07",X"8E",X"F8",X"07",X"48",
		X"A9",X"08",X"70",X"67",X"90",X"4D",X"B0",X"55",X"29",X"01",X"09",X"F0",X"9D",X"38",X"06",X"A9",
		X"02",X"D0",X"40",X"29",X"0F",X"09",X"90",X"D0",X"35",X"FF",X"FF",X"B9",X"83",X"C0",X"29",X"FB",
		X"99",X"83",X"C0",X"A9",X"3E",X"99",X"82",X"C0",X"B9",X"83",X"C0",X"09",X"04",X"99",X"83",X"C0",
		X"B9",X"82",X"C0",X"29",X"C1",X"1D",X"B8",X"05",X"99",X"82",X"C0",X"68",X"F0",X"0A",X"6A",X"90",
		X"75",X"68",X"AA",X"68",X"A8",X"68",X"28",X"60",X"18",X"60",X"29",X"01",X"09",X"60",X"9D",X"38",
		X"06",X"A9",X"0E",X"9D",X"B8",X"05",X"A9",X"01",X"48",X"D0",X"C0",X"A9",X"0C",X"9D",X"B8",X"05",
		X"A9",X"02",X"D0",X"F4",X"A9",X"30",X"9D",X"38",X"06",X"A9",X"06",X"9D",X"B8",X"05",X"A9",X"00",
		X"48",X"F0",X"A8",X"C9",X"10",X"B0",X"D2",X"9D",X"38",X"07",X"90",X"EA",X"A9",X"04",X"D0",X"EB",
		X"A9",X"40",X"D0",X"CA",X"A4",X"06",X"A9",X"60",X"85",X"06",X"20",X"06",X"00",X"84",X"06",X"BA",
		X"BD",X"00",X"01",X"AA",X"0A",X"0A",X"0A",X"0A",X"A8",X"A9",X"20",X"D0",X"C9",X"A9",X"70",X"D0",
		X"C5",X"48",X"A9",X"A0",X"D0",X"A8",X"29",X"0F",X"09",X"B0",X"D0",X"BA",X"A9",X"C0",X"D0",X"B6",
		X"A9",X"02",X"D0",X"B7",X"A2",X"03",X"38",X"60",X"FF",X"FF",X"FF",X"D6",X"FF",X"FF",X"FF",X"01",
		X"98",X"48",X"A5",X"06",X"48",X"A5",X"07",X"48",X"86",X"07",X"A9",X"27",X"85",X"06",X"20",X"58",
		X"FC",X"A0",X"00",X"B1",X"06",X"F0",X"06",X"20",X"ED",X"FD",X"C8",X"D0",X"F6",X"68",X"85",X"07",
		X"68",X"85",X"06",X"68",X"A8",X"D0",X"5B",X"C1",X"F0",X"F0",X"EC",X"E5",X"CD",X"EF",X"F5",X"F3",
		X"E5",X"8D",X"C3",X"EF",X"F0",X"F9",X"F2",X"E9",X"E7",X"E8",X"F4",X"A0",X"B1",X"B9",X"B8",X"B3",
		X"A0",X"E2",X"F9",X"A0",X"C1",X"F0",X"F0",X"EC",X"E5",X"A0",X"C3",X"EF",X"ED",X"F0",X"F5",X"F4",
		X"E5",X"F2",X"AC",X"A0",X"C9",X"EE",X"E3",X"AE",X"8D",X"8D",X"C2",X"E1",X"E3",X"E8",X"ED",X"E1",
		X"EE",X"AF",X"CD",X"E1",X"F2",X"EB",X"F3",X"AF",X"CD",X"E1",X"E3",X"CB",X"E1",X"F9",X"8D",X"00",
		X"B9",X"82",X"C0",X"29",X"F1",X"1D",X"B8",X"05",X"99",X"82",X"C0",X"68",X"30",X"0C",X"F0",X"80",
		X"D0",X"09",X"A9",X"00",X"9D",X"B8",X"05",X"48",X"F0",X"E6",X"60",X"BD",X"38",X"07",X"29",X"0F",
		X"09",X"20",X"9D",X"38",X"07",X"8A",X"48",X"48",X"48",X"48",X"A9",X"AA",X"48",X"BD",X"38",X"06",
		X"48",X"A9",X"0C",X"9D",X"B8",X"05",X"A9",X"00",X"48",X"F0",X"C5",X"A9",X"B3",X"48",X"AD",X"78",
		X"04",X"18",X"90",X"EC",X"A9",X"BC",X"48",X"AD",X"F8",X"04",X"18",X"90",X"E3",X"A9",X"81",X"48",
		X"7E",X"38",X"06",X"90",X"05",X"AD",X"78",X"05",X"B0",X"D6",X"8A",X"48",X"A9",X"D8",X"48",X"A9",
		X"0C",X"9D",X"B8",X"05",X"A9",X"01",X"48",X"D0",X"97",X"BD",X"38",X"06",X"8D",X"78",X"05",X"60",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"C2",
		X"BD",X"38",X"07",X"29",X"0F",X"09",X"40",X"9D",X"38",X"07",X"8A",X"48",X"48",X"48",X"A9",X"11",
		X"D0",X"27",X"A9",X"1E",X"48",X"A9",X"0C",X"9D",X"B8",X"05",X"A9",X"01",X"48",X"D0",X"51",X"AD",
		X"B3",X"FB",X"C9",X"06",X"D0",X"21",X"AD",X"19",X"C0",X"30",X"FB",X"AD",X"19",X"C0",X"10",X"FB",
		X"AD",X"19",X"C0",X"30",X"FB",X"A9",X"7F",X"D0",X"00",X"48",X"A9",X"50",X"48",X"A9",X"0C",X"9D",
		X"B8",X"05",X"A9",X"00",X"48",X"F0",X"29",X"A5",X"06",X"48",X"A5",X"07",X"48",X"98",X"48",X"A9",
		X"20",X"85",X"07",X"A0",X"00",X"84",X"06",X"A9",X"00",X"91",X"06",X"C8",X"D0",X"FB",X"E6",X"07",
		X"A5",X"07",X"C9",X"40",X"D0",X"F1",X"68",X"A8",X"A5",X"08",X"48",X"A9",X"00",X"F0",X"1C",X"FF",
		X"B9",X"82",X"C0",X"29",X"F1",X"1D",X"B8",X"05",X"99",X"82",X"C0",X"68",X"30",X"0A",X"F0",X"80",
		X"A9",X"00",X"9D",X"B8",X"05",X"48",X"F0",X"E8",X"60",X"D0",X"AE",X"A9",X"01",X"8D",X"D0",X"3F",
		X"8D",X"E0",X"3F",X"AD",X"57",X"C0",X"AD",X"54",X"C0",X"AD",X"52",X"C0",X"AD",X"50",X"C0",X"EA",
		X"85",X"06",X"85",X"07",X"85",X"08",X"E6",X"06",X"D0",X"0E",X"E6",X"07",X"D0",X"0C",X"E6",X"08",
		X"A5",X"08",X"C9",X"01",X"90",X"0A",X"B0",X"1F",X"08",X"28",X"08",X"28",X"A9",X"00",X"A5",X"00",
		X"AD",X"FF",X"CF",X"B9",X"82",X"C0",X"4A",X"EA",X"EA",X"B0",X"DB",X"AD",X"FF",X"CF",X"B9",X"82",
		X"C0",X"4A",X"A5",X"00",X"EA",X"B0",X"CF",X"68",X"85",X"08",X"68",X"85",X"07",X"68",X"85",X"06",
		X"A9",X"E3",X"D0",X"A5",X"AD",X"51",X"C0",X"AD",X"56",X"C0",X"18",X"90",X"93",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"C1",
		X"BD",X"38",X"06",X"C9",X"20",X"D0",X"06",X"A9",X"7F",X"69",X"01",X"70",X"01",X"B8",X"B9",X"82",
		X"C0",X"30",X"FB",X"B9",X"81",X"C0",X"29",X"FB",X"99",X"81",X"C0",X"A9",X"FF",X"99",X"80",X"C0",
		X"B9",X"81",X"C0",X"09",X"04",X"99",X"81",X"C0",X"BD",X"38",X"06",X"99",X"80",X"C0",X"B9",X"82",
		X"C0",X"09",X"20",X"99",X"82",X"C0",X"B9",X"82",X"C0",X"10",X"FB",X"29",X"DF",X"99",X"82",X"C0",
		X"70",X"44",X"BD",X"38",X"06",X"C9",X"30",X"D0",X"35",X"A9",X"00",X"9D",X"B8",X"04",X"9D",X"B8",
		X"03",X"9D",X"38",X"05",X"9D",X"38",X"04",X"F0",X"25",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"B9",X"82",X"C0",X"29",X"F1",X"1D",X"B8",X"05",X"99",X"82",X"C0",X"68",X"F0",X"82",X"A9",X"00",
		X"9D",X"B8",X"05",X"48",X"F0",X"EA",X"B9",X"81",X"C0",X"29",X"FB",X"99",X"81",X"C0",X"A9",X"00",
		X"99",X"80",X"C0",X"B9",X"81",X"C0",X"09",X"04",X"99",X"81",X"C0",X"B9",X"82",X"C0",X"0A",X"10",
		X"FA",X"B9",X"80",X"C0",X"9D",X"38",X"06",X"B9",X"82",X"C0",X"09",X"10",X"99",X"82",X"C0",X"B9",
		X"82",X"C0",X"0A",X"30",X"FA",X"B9",X"82",X"C0",X"29",X"EF",X"99",X"82",X"C0",X"BD",X"B8",X"06",
		X"29",X"F1",X"1D",X"38",X"06",X"9D",X"B8",X"06",X"29",X"0E",X"D0",X"B2",X"A9",X"00",X"9D",X"B8",
		X"05",X"A9",X"02",X"48",X"D0",X"9A",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"C3",
		X"E4",X"37",X"D0",X"2D",X"A9",X"07",X"C5",X"36",X"F0",X"27",X"85",X"36",X"68",X"C9",X"8D",X"F0",
		X"74",X"29",X"01",X"09",X"80",X"9D",X"38",X"07",X"8A",X"48",X"A9",X"84",X"48",X"BD",X"38",X"07",
		X"4A",X"A9",X"80",X"B0",X"01",X"0A",X"48",X"A9",X"0C",X"9D",X"B8",X"05",X"A9",X"00",X"48",X"F0",
		X"3F",X"E4",X"39",X"D0",X"D7",X"A9",X"05",X"85",X"38",X"BD",X"38",X"07",X"29",X"01",X"D0",X"14",
		X"68",X"68",X"68",X"68",X"A9",X"00",X"9D",X"B8",X"03",X"9D",X"B8",X"04",X"9D",X"38",X"04",X"9D",
		X"38",X"05",X"F0",X"3C",X"BD",X"38",X"07",X"29",X"01",X"09",X"80",X"9D",X"38",X"07",X"8A",X"48",
		X"A9",X"A1",X"48",X"A9",X"10",X"48",X"A9",X"0C",X"D0",X"30",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"B9",X"82",X"C0",X"29",X"F1",X"1D",X"B8",X"05",X"99",X"82",X"C0",X"68",X"30",X"11",X"F0",X"80",
		X"6A",X"B0",X"89",X"90",X"B4",X"A9",X"00",X"9D",X"B8",X"05",X"A9",X"01",X"48",X"D0",X"E1",X"60",
		X"A9",X"C0",X"9D",X"B8",X"06",X"8C",X"22",X"02",X"A9",X"0A",X"9D",X"B8",X"05",X"A9",X"00",X"48",
		X"F0",X"CE",X"68",X"68",X"68",X"68",X"A9",X"05",X"9D",X"38",X"06",X"B9",X"81",X"C0",X"29",X"FB",
		X"99",X"81",X"C0",X"A9",X"00",X"99",X"80",X"C0",X"B9",X"81",X"C0",X"09",X"04",X"99",X"81",X"C0",
		X"B9",X"82",X"C0",X"0A",X"10",X"FA",X"B9",X"80",X"C0",X"48",X"B9",X"82",X"C0",X"09",X"10",X"99",
		X"82",X"C0",X"B9",X"82",X"C0",X"0A",X"30",X"FA",X"B9",X"82",X"C0",X"29",X"EF",X"99",X"82",X"C0",
		X"DE",X"38",X"06",X"D0",X"DB",X"68",X"9D",X"B8",X"06",X"68",X"9D",X"38",X"05",X"68",X"9D",X"38",
		X"04",X"68",X"9D",X"B8",X"04",X"68",X"9D",X"B8",X"03",X"18",X"90",X"99",X"FF",X"FF",X"FF",X"C8",
		X"8A",X"48",X"48",X"48",X"A9",X"12",X"48",X"BC",X"B8",X"03",X"BD",X"B8",X"04",X"AA",X"98",X"A0",
		X"05",X"D0",X"6D",X"AE",X"F8",X"07",X"A9",X"24",X"48",X"BC",X"38",X"04",X"BD",X"38",X"05",X"AA",
		X"98",X"A0",X"0C",X"D0",X"5B",X"AE",X"F8",X"07",X"A9",X"43",X"48",X"AD",X"00",X"C0",X"0A",X"08",
		X"BD",X"B8",X"06",X"2A",X"2A",X"2A",X"29",X"03",X"49",X"03",X"38",X"69",X"00",X"28",X"A2",X"00",
		X"A0",X"10",X"D0",X"4D",X"A9",X"8D",X"8D",X"11",X"02",X"48",X"A9",X"11",X"48",X"48",X"A9",X"00",
		X"F0",X"12",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"AE",X"F8",X"07",X"AC",X"22",X"02",X"9D",X"B8",X"05",X"A9",X"01",X"48",
		X"B9",X"82",X"C0",X"29",X"F1",X"1D",X"B8",X"05",X"99",X"82",X"C0",X"68",X"30",X"4E",X"F0",X"80",
		X"E0",X"80",X"90",X"0D",X"49",X"FF",X"69",X"00",X"48",X"8A",X"49",X"FF",X"69",X"00",X"AA",X"68",
		X"38",X"8D",X"21",X"02",X"8E",X"20",X"02",X"A9",X"AB",X"90",X"02",X"A9",X"AD",X"48",X"A9",X"AC",
		X"99",X"01",X"02",X"A2",X"11",X"A9",X"00",X"18",X"2A",X"C9",X"0A",X"90",X"02",X"E9",X"0A",X"2E",
		X"21",X"02",X"2E",X"20",X"02",X"CA",X"D0",X"F0",X"09",X"B0",X"99",X"00",X"02",X"88",X"F0",X"08",
		X"C0",X"07",X"F0",X"04",X"C0",X"0E",X"D0",X"DB",X"68",X"99",X"00",X"02",X"60",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"CD",
		X"B8",X"50",X"13",X"BD",X"38",X"07",X"29",X"01",X"F0",X"47",X"A9",X"10",X"48",X"A9",X"05",X"9D",
		X"38",X"06",X"A9",X"7F",X"69",X"01",X"B9",X"82",X"C0",X"30",X"FB",X"B9",X"81",X"C0",X"29",X"FB",
		X"99",X"81",X"C0",X"A9",X"FF",X"99",X"80",X"C0",X"B9",X"81",X"C0",X"09",X"04",X"99",X"81",X"C0",
		X"68",X"99",X"80",X"C0",X"B9",X"82",X"C0",X"09",X"20",X"99",X"82",X"C0",X"B9",X"82",X"C0",X"10",
		X"FB",X"29",X"DF",X"99",X"82",X"C0",X"70",X"3F",X"70",X"07",X"BD",X"38",X"07",X"4A",X"4A",X"4A",
		X"4A",X"B8",X"9D",X"B8",X"05",X"F0",X"02",X"A9",X"80",X"48",X"50",X"14",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"B9",X"82",X"C0",X"29",X"F1",X"1D",X"B8",X"05",X"99",X"82",X"C0",X"68",X"F0",X"82",X"C9",X"02",
		X"F0",X"81",X"D0",X"02",X"F0",X"C2",X"B8",X"B9",X"81",X"C0",X"29",X"FB",X"99",X"81",X"C0",X"A9",
		X"00",X"99",X"80",X"C0",X"B9",X"81",X"C0",X"09",X"04",X"99",X"81",X"C0",X"B9",X"82",X"C0",X"0A",
		X"10",X"FA",X"B9",X"80",X"C0",X"70",X"05",X"9D",X"38",X"06",X"50",X"01",X"48",X"B9",X"82",X"C0",
		X"09",X"10",X"99",X"82",X"C0",X"B9",X"82",X"C0",X"0A",X"30",X"FA",X"B9",X"82",X"C0",X"29",X"EF",
		X"99",X"82",X"C0",X"50",X"19",X"DE",X"38",X"06",X"D0",X"D2",X"68",X"9D",X"B8",X"06",X"68",X"9D",
		X"38",X"05",X"68",X"9D",X"38",X"04",X"68",X"9D",X"B8",X"04",X"68",X"9D",X"B8",X"03",X"A9",X"00",
		X"F0",X"A2",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"C1",
		X"BD",X"38",X"06",X"C9",X"40",X"F0",X"22",X"C9",X"60",X"F0",X"0D",X"C9",X"61",X"F0",X"09",X"C9",
		X"A0",X"D0",X"2E",X"48",X"A9",X"02",X"D0",X"45",X"AD",X"F8",X"05",X"48",X"AD",X"78",X"05",X"48",
		X"AD",X"F8",X"04",X"48",X"AD",X"78",X"04",X"B0",X"0F",X"BD",X"38",X"05",X"48",X"BD",X"38",X"04",
		X"48",X"BD",X"B8",X"04",X"48",X"BD",X"B8",X"03",X"48",X"BD",X"38",X"06",X"48",X"A9",X"05",X"D0",
		X"1C",X"29",X"0C",X"4A",X"4A",X"4A",X"B0",X"3E",X"4A",X"90",X"0C",X"AD",X"78",X"05",X"48",X"BD",
		X"38",X"06",X"48",X"A9",X"02",X"D0",X"06",X"BD",X"38",X"06",X"48",X"A9",X"01",X"9D",X"38",X"06",
		X"D0",X"4F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"B9",X"82",X"C0",X"29",X"F1",X"1D",X"B8",X"05",X"99",X"82",X"C0",X"68",X"D0",X"82",X"A9",X"00",
		X"9D",X"B8",X"05",X"48",X"F0",X"EA",X"4A",X"B0",X"13",X"AD",X"F8",X"04",X"48",X"AD",X"78",X"04",
		X"48",X"BD",X"38",X"06",X"48",X"A9",X"03",X"9D",X"38",X"06",X"D0",X"15",X"AD",X"78",X"05",X"48",
		X"AD",X"F8",X"04",X"48",X"AD",X"78",X"04",X"48",X"BD",X"38",X"06",X"48",X"A9",X"04",X"9D",X"38",
		X"06",X"B9",X"82",X"C0",X"30",X"FB",X"B9",X"81",X"C0",X"29",X"FB",X"99",X"81",X"C0",X"A9",X"FF",
		X"99",X"80",X"C0",X"B9",X"81",X"C0",X"09",X"04",X"99",X"81",X"C0",X"68",X"99",X"80",X"C0",X"B9",
		X"82",X"C0",X"09",X"20",X"99",X"82",X"C0",X"B9",X"82",X"C0",X"10",X"FB",X"29",X"DF",X"99",X"82",
		X"C0",X"DE",X"38",X"06",X"F0",X"98",X"B9",X"82",X"C0",X"30",X"FB",X"10",X"D6",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"CE");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
