library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity applemouse_mcu_rom is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(10 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of applemouse_mcu_rom is
	type rom is array(0 to  2047) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"03",X"02",X"FD",X"B6",X"00",X"16",X"02",X"02",X"02",X"FD",X"17",X"02",X"81",X"00",X"02",X"FD",
		X"B7",X"00",X"14",X"02",X"01",X"02",X"FD",X"15",X"02",X"81",X"02",X"08",X"01",X"04",X"CC",X"04",
		X"6C",X"00",X"CC",X"04",X"73",X"00",X"CC",X"04",X"DC",X"00",X"CC",X"05",X"1B",X"00",X"CC",X"05",
		X"2C",X"00",X"CC",X"05",X"47",X"00",X"CC",X"05",X"74",X"00",X"CC",X"05",X"90",X"00",X"CC",X"05",
		X"A7",X"00",X"CC",X"05",X"B0",X"00",X"CC",X"06",X"17",X"00",X"CC",X"06",X"1F",X"00",X"CC",X"06",
		X"26",X"00",X"CC",X"06",X"7A",X"00",X"CC",X"06",X"7A",X"00",X"CC",X"06",X"48",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"A6",X"00",X"B7",X"00",X"B7",X"02",X"B7",X"04",X"A6",X"0C",X"B7",X"06",X"A6",X"40",X"B7",X"01",
		X"B7",X"05",X"C6",X"06",X"C7",X"B7",X"51",X"C6",X"06",X"C9",X"B7",X"50",X"C6",X"06",X"C3",X"B7",
		X"53",X"C6",X"06",X"C5",X"B7",X"52",X"A6",X"01",X"B7",X"57",X"A6",X"00",X"B7",X"54",X"B7",X"55",
		X"CC",X"04",X"F9",X"03",X"02",X"0D",X"CD",X"00",X"83",X"B7",X"59",X"44",X"44",X"A4",X"3C",X"97",
		X"DC",X"00",X"9E",X"B6",X"01",X"A4",X"0F",X"B8",X"44",X"27",X"E8",X"01",X"58",X"5B",X"B7",X"45",
		X"B8",X"44",X"B7",X"44",X"01",X"5D",X"08",X"A4",X"0A",X"B4",X"45",X"27",X"4C",X"B7",X"45",X"A6",
		X"20",X"B7",X"5A",X"A6",X"02",X"B7",X"5B",X"AE",X"01",X"B6",X"45",X"D4",X"00",X"9A",X"27",X"36",
		X"B6",X"44",X"D4",X"00",X"9C",X"27",X"18",X"E6",X"42",X"E1",X"4D",X"26",X"09",X"E6",X"40",X"E1",
		X"4B",X"26",X"03",X"CC",X"04",X"4C",X"6C",X"42",X"26",X"02",X"6C",X"40",X"CC",X"04",X"66",X"E6",
		X"42",X"E1",X"49",X"26",X"09",X"E6",X"40",X"E1",X"47",X"26",X"03",X"CC",X"04",X"66",X"E6",X"42",
		X"26",X"02",X"6A",X"40",X"6A",X"42",X"5A",X"27",X"C0",X"CC",X"03",X"F3",X"B6",X"59",X"B7",X"58",
		X"CC",X"04",X"03",X"A6",X"FF",X"B7",X"04",X"B6",X"42",X"00",X"02",X"FD",X"B7",X"00",X"14",X"02",
		X"01",X"02",X"FD",X"15",X"02",X"B6",X"40",X"00",X"02",X"FD",X"B7",X"00",X"14",X"02",X"01",X"02",
		X"FD",X"15",X"02",X"B6",X"43",X"00",X"02",X"FD",X"B7",X"00",X"14",X"02",X"01",X"02",X"FD",X"15",
		X"02",X"B6",X"41",X"00",X"02",X"FD",X"B7",X"00",X"14",X"02",X"01",X"02",X"FD",X"15",X"02",X"B6",
		X"01",X"A8",X"80",X"48",X"36",X"46",X"B6",X"46",X"A4",X"C0",X"BA",X"5A",X"00",X"02",X"FD",X"B7",
		X"00",X"14",X"02",X"01",X"02",X"FD",X"15",X"02",X"A6",X"00",X"B7",X"5A",X"B7",X"04",X"03",X"5D",
		X"08",X"B7",X"40",X"B7",X"42",X"B7",X"41",X"B7",X"43",X"CC",X"04",X"03",X"1C",X"01",X"A6",X"FF",
		X"B7",X"04",X"B6",X"5C",X"00",X"02",X"FD",X"B7",X"00",X"14",X"02",X"01",X"02",X"FD",X"15",X"02",
		X"A6",X"00",X"B7",X"5C",X"B7",X"04",X"CC",X"04",X"03",X"B7",X"5B",X"B7",X"5C",X"B7",X"58",X"B7",
		X"5D",X"B7",X"47",X"B7",X"49",X"B7",X"48",X"B7",X"4A",X"A6",X"03",X"B7",X"4B",X"B7",X"4C",X"A6",
		X"FF",X"B7",X"4D",X"B7",X"4E",X"B6",X"01",X"A4",X"0F",X"B7",X"44",X"A6",X"00",X"B7",X"46",X"B7",
		X"5A",X"B7",X"40",X"B7",X"42",X"B7",X"41",X"B7",X"43",X"CC",X"04",X"03",X"CD",X"00",X"80",X"B7",
		X"42",X"CD",X"00",X"80",X"B7",X"40",X"CD",X"00",X"80",X"B7",X"43",X"CD",X"00",X"80",X"B7",X"41",
		X"A6",X"00",X"B7",X"5A",X"CC",X"04",X"03",X"9B",X"1D",X"09",X"B6",X"57",X"B7",X"56",X"B6",X"53",
		X"4C",X"B7",X"4F",X"A6",X"00",X"B7",X"5B",X"B7",X"5C",X"1C",X"01",X"CD",X"00",X"8D",X"03",X"02",
		X"FD",X"A6",X"FF",X"B7",X"08",X"1F",X"09",X"9A",X"B6",X"52",X"B7",X"08",X"CD",X"00",X"83",X"A6",
		X"00",X"CC",X"04",X"FD",X"B6",X"59",X"A4",X"01",X"97",X"CD",X"00",X"80",X"E7",X"49",X"CD",X"00",
		X"80",X"E7",X"4D",X"CD",X"00",X"80",X"E7",X"47",X"CD",X"00",X"80",X"E7",X"4B",X"CC",X"04",X"03",
		X"B6",X"49",X"B7",X"42",X"B6",X"47",X"B7",X"40",X"B6",X"4A",X"B7",X"43",X"B6",X"48",X"B7",X"41",
		X"A6",X"00",X"B7",X"5A",X"CC",X"04",X"03",X"A6",X"01",X"B7",X"58",X"A6",X"00",X"CC",X"04",X"FF",
		X"1C",X"09",X"B6",X"59",X"A4",X"01",X"97",X"D6",X"06",X"C5",X"B7",X"52",X"D6",X"06",X"C3",X"B7",
		X"53",X"D6",X"06",X"C9",X"B7",X"50",X"D6",X"06",X"C7",X"B7",X"51",X"B6",X"59",X"A4",X"04",X"27",
		X"18",X"CD",X"00",X"80",X"B7",X"54",X"CD",X"00",X"80",X"B7",X"55",X"B6",X"52",X"BB",X"54",X"B7",
		X"52",X"B6",X"53",X"B9",X"55",X"B7",X"53",X"20",X"06",X"A6",X"00",X"B7",X"54",X"B7",X"55",X"B6",
		X"59",X"A4",X"02",X"27",X"0E",X"B6",X"52",X"CB",X"06",X"C2",X"B7",X"52",X"B6",X"53",X"C9",X"06",
		X"C1",X"B7",X"53",X"B6",X"59",X"A4",X"08",X"27",X"07",X"CD",X"00",X"80",X"B7",X"57",X"20",X"04",
		X"A6",X"01",X"B7",X"57",X"CC",X"04",X"03",X"CD",X"00",X"80",X"B7",X"57",X"CC",X"04",X"03",X"B6",
		X"59",X"B7",X"5D",X"CC",X"04",X"03",X"9B",X"1D",X"09",X"A6",X"00",X"B7",X"5B",X"B7",X"5C",X"1C",
		X"01",X"B6",X"57",X"B7",X"56",X"B6",X"55",X"4C",X"B7",X"08",X"A6",X"FF",X"B7",X"08",X"1F",X"09",
		X"9A",X"B6",X"54",X"B7",X"08",X"CC",X"04",X"03",X"CD",X"00",X"80",X"B7",X"60",X"CD",X"00",X"80",
		X"B7",X"5F",X"A6",X"81",X"B7",X"61",X"B6",X"59",X"A4",X"01",X"26",X"12",X"A6",X"FF",X"B7",X"04",
		X"A6",X"C6",X"B7",X"5E",X"BD",X"5E",X"CD",X"00",X"8D",X"3F",X"04",X"CC",X"04",X"03",X"A6",X"C7",
		X"B7",X"5E",X"CD",X"00",X"80",X"BD",X"5E",X"CC",X"04",X"03",X"CC",X"04",X"03",X"1F",X"09",X"3A",
		X"4F",X"26",X"3C",X"B6",X"08",X"B0",X"50",X"B7",X"08",X"B6",X"4F",X"B2",X"51",X"4C",X"B7",X"4F",
		X"3A",X"56",X"26",X"2B",X"B6",X"57",X"B7",X"56",X"B6",X"01",X"2B",X"04",X"A6",X"0C",X"20",X"04",
		X"A6",X"08",X"20",X"00",X"BA",X"5B",X"00",X"58",X"04",X"A4",X"08",X"20",X"04",X"A4",X"0E",X"20",
		X"00",X"B4",X"58",X"27",X"02",X"1D",X"01",X"BA",X"5C",X"B7",X"5C",X"A6",X"00",X"B7",X"5B",X"80",
		X"80",X"FC",X"8E",X"41",X"4E",X"A2",X"4E",X"DF",X"D9",X"C7",X"6E",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"41",X"50",X"50",X"4C",X"45",X"4D",X"4F",X"55",X"53",
		X"45",X"8D",X"43",X"4F",X"50",X"59",X"52",X"49",X"47",X"48",X"54",X"20",X"31",X"39",X"38",X"33",
		X"20",X"42",X"59",X"20",X"41",X"50",X"50",X"4C",X"45",X"20",X"43",X"4F",X"4D",X"50",X"55",X"54",
		X"45",X"52",X"2C",X"20",X"49",X"4E",X"43",X"2E",X"8D",X"41",X"4C",X"4C",X"20",X"52",X"49",X"47",
		X"48",X"54",X"53",X"20",X"52",X"45",X"53",X"45",X"52",X"56",X"45",X"44",X"8D",X"4D",X"41",X"52",
		X"4B",X"53",X"2F",X"4D",X"41",X"43",X"44",X"4F",X"55",X"47",X"41",X"4C",X"4C",X"2F",X"4D",X"41",
		X"43",X"4B",X"41",X"59",X"2F",X"42",X"41",X"43",X"48",X"4D",X"41",X"4E",X"8D",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"06",X"7D",X"06",X"C0",X"06",X"C0",X"03",X"C0");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
