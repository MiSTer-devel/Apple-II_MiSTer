library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity main_roms is
 port (
   addr : in  unsigned(13 downto 0);
   clk  : in  std_logic;
   dout : out unsigned(7 downto 0));
end main_roms;

architecture rtl of main_roms is
  type rom_array is array(0 to 12287) of unsigned(7 downto 0);

  constant ROM : rom_array := (
     X"6f", X"d8", X"65", X"d7", X"f8", X"dc", X"94", X"d9",
     X"b1", X"db", X"30", X"f3", X"d8", X"df", X"e1", X"db",
     X"8f", X"f3", X"98", X"f3", X"e4", X"f1", X"dd", X"f1",
     X"d4", X"f1", X"24", X"f2", X"31", X"f2", X"40", X"f2",
     X"d7", X"f3", X"e1", X"f3", X"e8", X"f6", X"fd", X"f6",
     X"68", X"f7", X"6e", X"f7", X"e6", X"f7", X"57", X"fc",
     X"20", X"f7", X"26", X"f7", X"74", X"f7", X"6c", X"f2",
     X"6e", X"f2", X"72", X"f2", X"76", X"f2", X"7f", X"f2",
     X"4e", X"f2", X"6a", X"d9", X"55", X"f2", X"85", X"f2",
     X"a5", X"f2", X"ca", X"f2", X"17", X"f3", X"bb", X"f3",
     X"9e", X"f3", X"61", X"f2", X"45", X"da", X"3d", X"d9",
     X"11", X"d9", X"c8", X"d9", X"48", X"d8", X"f4", X"03",
     X"20", X"d9", X"6a", X"d9", X"db", X"d9", X"6d", X"d8",
     X"eb", X"d9", X"83", X"e7", X"c8", X"d8", X"af", X"d8",
     X"12", X"e3", X"7a", X"e7", X"d4", X"da", X"95", X"d8",
     X"a4", X"d6", X"69", X"d6", X"9f", X"db", X"48", X"d6",
     X"90", X"eb", X"23", X"ec", X"af", X"eb", X"0a", X"00",
     X"de", X"e2", X"12", X"d4", X"cd", X"df", X"ff", X"e2",
     X"8d", X"ee", X"ae", X"ef", X"41", X"e9", X"09", X"ef",
     X"ea", X"ef", X"f1", X"ef", X"3a", X"f0", X"9e", X"f0",
     X"64", X"e7", X"d6", X"e6", X"c5", X"e3", X"07", X"e7",
     X"e5", X"e6", X"46", X"e6", X"5a", X"e6", X"86", X"e6",
     X"91", X"e6", X"79", X"c0", X"e7", X"79", X"a9", X"e7",
     X"7b", X"81", X"e9", X"7b", X"68", X"ea", X"7d", X"96",
     X"ee", X"50", X"54", X"df", X"46", X"4e", X"df", X"7f",
     X"cf", X"ee", X"7f", X"97", X"de", X"64", X"64", X"df",
     X"45", X"4e", X"c4", X"46", X"4f", X"d2", X"4e", X"45",
     X"58", X"d4", X"44", X"41", X"54", X"c1", X"49", X"4e",
     X"50", X"55", X"d4", X"44", X"45", X"cc", X"44", X"49",
     X"cd", X"52", X"45", X"41", X"c4", X"47", X"d2", X"54",
     X"45", X"58", X"d4", X"50", X"52", X"a3", X"49", X"4e",
     X"a3", X"43", X"41", X"4c", X"cc", X"50", X"4c", X"4f",
     X"d4", X"48", X"4c", X"49", X"ce", X"56", X"4c", X"49",
     X"ce", X"48", X"47", X"52", X"b2", X"48", X"47", X"d2",
     X"48", X"43", X"4f", X"4c", X"4f", X"52", X"bd", X"48",
     X"50", X"4c", X"4f", X"d4", X"44", X"52", X"41", X"d7",
     X"58", X"44", X"52", X"41", X"d7", X"48", X"54", X"41",
     X"c2", X"48", X"4f", X"4d", X"c5", X"52", X"4f", X"54",
     X"bd", X"53", X"43", X"41", X"4c", X"45", X"bd", X"53",
     X"48", X"4c", X"4f", X"41", X"c4", X"54", X"52", X"41",
     X"43", X"c5", X"4e", X"4f", X"54", X"52", X"41", X"43",
     X"c5", X"4e", X"4f", X"52", X"4d", X"41", X"cc", X"49",
     X"4e", X"56", X"45", X"52", X"53", X"c5", X"46", X"4c",
     X"41", X"53", X"c8", X"43", X"4f", X"4c", X"4f", X"52",
     X"bd", X"50", X"4f", X"d0", X"56", X"54", X"41", X"c2",
     X"48", X"49", X"4d", X"45", X"4d", X"ba", X"4c", X"4f",
     X"4d", X"45", X"4d", X"ba", X"4f", X"4e", X"45", X"52",
     X"d2", X"52", X"45", X"53", X"55", X"4d", X"c5", X"52",
     X"45", X"43", X"41", X"4c", X"cc", X"53", X"54", X"4f",
     X"52", X"c5", X"53", X"50", X"45", X"45", X"44", X"bd",
     X"4c", X"45", X"d4", X"47", X"4f", X"54", X"cf", X"52",
     X"55", X"ce", X"49", X"c6", X"52", X"45", X"53", X"54",
     X"4f", X"52", X"c5", X"a6", X"47", X"4f", X"53", X"55",
     X"c2", X"52", X"45", X"54", X"55", X"52", X"ce", X"52",
     X"45", X"cd", X"53", X"54", X"4f", X"d0", X"4f", X"ce",
     X"57", X"41", X"49", X"d4", X"4c", X"4f", X"41", X"c4",
     X"53", X"41", X"56", X"c5", X"44", X"45", X"c6", X"50",
     X"4f", X"4b", X"c5", X"50", X"52", X"49", X"4e", X"d4",
     X"43", X"4f", X"4e", X"d4", X"4c", X"49", X"53", X"d4",
     X"43", X"4c", X"45", X"41", X"d2", X"47", X"45", X"d4",
     X"4e", X"45", X"d7", X"54", X"41", X"42", X"a8", X"54",
     X"cf", X"46", X"ce", X"53", X"50", X"43", X"a8", X"54",
     X"48", X"45", X"ce", X"41", X"d4", X"4e", X"4f", X"d4",
     X"53", X"54", X"45", X"d0", X"ab", X"ad", X"aa", X"af",
     X"de", X"41", X"4e", X"c4", X"4f", X"d2", X"be", X"bd",
     X"bc", X"53", X"47", X"ce", X"49", X"4e", X"d4", X"41",
     X"42", X"d3", X"55", X"53", X"d2", X"46", X"52", X"c5",
     X"53", X"43", X"52", X"4e", X"a8", X"50", X"44", X"cc",
     X"50", X"4f", X"d3", X"53", X"51", X"d2", X"52", X"4e",
     X"c4", X"4c", X"4f", X"c7", X"45", X"58", X"d0", X"43",
     X"4f", X"d3", X"53", X"49", X"ce", X"54", X"41", X"ce",
     X"41", X"54", X"ce", X"50", X"45", X"45", X"cb", X"4c",
     X"45", X"ce", X"53", X"54", X"52", X"a4", X"56", X"41",
     X"cc", X"41", X"53", X"c3", X"43", X"48", X"52", X"a4",
     X"4c", X"45", X"46", X"54", X"a4", X"52", X"49", X"47",
     X"48", X"54", X"a4", X"4d", X"49", X"44", X"a4", X"00",
     X"4e", X"45", X"58", X"54", X"20", X"57", X"49", X"54",
     X"48", X"4f", X"55", X"54", X"20", X"46", X"4f", X"d2",
     X"53", X"59", X"4e", X"54", X"41", X"d8", X"52", X"45",
     X"54", X"55", X"52", X"4e", X"20", X"57", X"49", X"54",
     X"48", X"4f", X"55", X"54", X"20", X"47", X"4f", X"53",
     X"55", X"c2", X"4f", X"55", X"54", X"20", X"4f", X"46",
     X"20", X"44", X"41", X"54", X"c1", X"49", X"4c", X"4c",
     X"45", X"47", X"41", X"4c", X"20", X"51", X"55", X"41",
     X"4e", X"54", X"49", X"54", X"d9", X"4f", X"56", X"45",
     X"52", X"46", X"4c", X"4f", X"d7", X"4f", X"55", X"54",
     X"20", X"4f", X"46", X"20", X"4d", X"45", X"4d", X"4f",
     X"52", X"d9", X"55", X"4e", X"44", X"45", X"46", X"27",
     X"44", X"20", X"53", X"54", X"41", X"54", X"45", X"4d",
     X"45", X"4e", X"d4", X"42", X"41", X"44", X"20", X"53",
     X"55", X"42", X"53", X"43", X"52", X"49", X"50", X"d4",
     X"52", X"45", X"44", X"49", X"4d", X"27", X"44", X"20",
     X"41", X"52", X"52", X"41", X"d9", X"44", X"49", X"56",
     X"49", X"53", X"49", X"4f", X"4e", X"20", X"42", X"59",
     X"20", X"5a", X"45", X"52", X"cf", X"49", X"4c", X"4c",
     X"45", X"47", X"41", X"4c", X"20", X"44", X"49", X"52",
     X"45", X"43", X"d4", X"54", X"59", X"50", X"45", X"20",
     X"4d", X"49", X"53", X"4d", X"41", X"54", X"43", X"c8",
     X"53", X"54", X"52", X"49", X"4e", X"47", X"20", X"54",
     X"4f", X"4f", X"20", X"4c", X"4f", X"4e", X"c7", X"46",
     X"4f", X"52", X"4d", X"55", X"4c", X"41", X"20", X"54",
     X"4f", X"4f", X"20", X"43", X"4f", X"4d", X"50", X"4c",
     X"45", X"d8", X"43", X"41", X"4e", X"27", X"54", X"20",
     X"43", X"4f", X"4e", X"54", X"49", X"4e", X"55", X"c5",
     X"55", X"4e", X"44", X"45", X"46", X"27", X"44", X"20",
     X"46", X"55", X"4e", X"43", X"54", X"49", X"4f", X"ce",
     X"20", X"45", X"52", X"52", X"4f", X"52", X"07", X"00",
     X"20", X"49", X"4e", X"20", X"00", X"0d", X"42", X"52",
     X"45", X"41", X"4b", X"07", X"00", X"ba", X"e8", X"e8",
     X"e8", X"e8", X"bd", X"01", X"01", X"c9", X"81", X"d0",
     X"21", X"a5", X"86", X"d0", X"0a", X"bd", X"02", X"01",
     X"85", X"85", X"bd", X"03", X"01", X"85", X"86", X"dd",
     X"03", X"01", X"d0", X"07", X"a5", X"85", X"dd", X"02",
     X"01", X"f0", X"07", X"8a", X"18", X"69", X"12", X"aa",
     X"d0", X"d8", X"60", X"20", X"e3", X"d3", X"85", X"6d",
     X"84", X"6e", X"38", X"a5", X"96", X"e5", X"9b", X"85",
     X"5e", X"a8", X"a5", X"97", X"e5", X"9c", X"aa", X"e8",
     X"98", X"f0", X"23", X"a5", X"96", X"38", X"e5", X"5e",
     X"85", X"96", X"b0", X"03", X"c6", X"97", X"38", X"a5",
     X"94", X"e5", X"5e", X"85", X"94", X"b0", X"08", X"c6",
     X"95", X"90", X"04", X"b1", X"96", X"91", X"94", X"88",
     X"d0", X"f9", X"b1", X"96", X"91", X"94", X"c6", X"97",
     X"c6", X"95", X"ca", X"d0", X"f2", X"60", X"0a", X"69",
     X"36", X"b0", X"35", X"85", X"5e", X"ba", X"e4", X"5e",
     X"90", X"2e", X"60", X"c4", X"70", X"90", X"28", X"d0",
     X"04", X"c5", X"6f", X"90", X"22", X"48", X"a2", X"09",
     X"98", X"48", X"b5", X"93", X"ca", X"10", X"fa", X"20",
     X"84", X"e4", X"a2", X"f7", X"68", X"95", X"9d", X"e8",
     X"30", X"fa", X"68", X"a8", X"68", X"c4", X"70", X"90",
     X"06", X"d0", X"05", X"c5", X"6f", X"b0", X"01", X"60",
     X"a2", X"4d", X"24", X"d8", X"10", X"03", X"4c", X"e9",
     X"f2", X"20", X"fb", X"da", X"20", X"5a", X"db", X"bd",
     X"60", X"d2", X"48", X"20", X"5c", X"db", X"e8", X"68",
     X"10", X"f5", X"20", X"83", X"d6", X"a9", X"50", X"a0",
     X"d3", X"20", X"3a", X"db", X"a4", X"76", X"c8", X"f0",
     X"03", X"20", X"19", X"ed", X"20", X"fb", X"da", X"a2",
     X"dd", X"20", X"2e", X"d5", X"86", X"b8", X"84", X"b9",
     X"46", X"d8", X"20", X"b1", X"00", X"aa", X"f0", X"ec",
     X"a2", X"ff", X"86", X"76", X"90", X"06", X"20", X"59",
     X"d5", X"4c", X"05", X"d8", X"a6", X"af", X"86", X"69",
     X"a6", X"b0", X"86", X"6a", X"20", X"0c", X"da", X"20",
     X"59", X"d5", X"84", X"0f", X"20", X"1a", X"d6", X"90",
     X"44", X"a0", X"01", X"b1", X"9b", X"85", X"5f", X"a5",
     X"69", X"85", X"5e", X"a5", X"9c", X"85", X"61", X"a5",
     X"9b", X"88", X"f1", X"9b", X"18", X"65", X"69", X"85",
     X"69", X"85", X"60", X"a5", X"6a", X"69", X"ff", X"85",
     X"6a", X"e5", X"9c", X"aa", X"38", X"a5", X"9b", X"e5",
     X"69", X"a8", X"b0", X"03", X"e8", X"c6", X"61", X"18",
     X"65", X"5e", X"90", X"03", X"c6", X"5f", X"18", X"b1",
     X"5e", X"91", X"60", X"c8", X"d0", X"f9", X"e6", X"5f",
     X"e6", X"61", X"ca", X"d0", X"f2", X"ad", X"00", X"02",
     X"f0", X"38", X"a5", X"73", X"a4", X"74", X"85", X"6f",
     X"84", X"70", X"a5", X"69", X"85", X"96", X"65", X"0f",
     X"85", X"94", X"a4", X"6a", X"84", X"97", X"90", X"01",
     X"c8", X"84", X"95", X"20", X"93", X"d3", X"a5", X"50",
     X"a4", X"51", X"8d", X"fe", X"01", X"8c", X"ff", X"01",
     X"a5", X"6d", X"a4", X"6e", X"85", X"69", X"84", X"6a",
     X"a4", X"0f", X"b9", X"fb", X"01", X"88", X"91", X"9b",
     X"d0", X"f8", X"20", X"65", X"d6", X"a5", X"67", X"a4",
     X"68", X"85", X"5e", X"84", X"5f", X"18", X"a0", X"01",
     X"b1", X"5e", X"d0", X"0b", X"a5", X"69", X"85", X"af",
     X"a5", X"6a", X"85", X"b0", X"4c", X"3c", X"d4", X"a0",
     X"04", X"c8", X"b1", X"5e", X"d0", X"fb", X"c8", X"98",
     X"65", X"5e", X"aa", X"a0", X"00", X"91", X"5e", X"a5",
     X"5f", X"69", X"00", X"c8", X"91", X"5e", X"86", X"5e",
     X"85", X"5f", X"90", X"d2", X"a2", X"80", X"86", X"33",
     X"20", X"6a", X"fd", X"e0", X"ef", X"90", X"02", X"a2",
     X"ef", X"a9", X"00", X"9d", X"00", X"02", X"8a", X"f0",
     X"0b", X"bd", X"ff", X"01", X"29", X"7f", X"9d", X"ff",
     X"01", X"ca", X"d0", X"f5", X"a9", X"00", X"a2", X"ff",
     X"a0", X"01", X"60", X"20", X"0c", X"fd", X"29", X"7f",
     X"60", X"a6", X"b8", X"ca", X"a0", X"04", X"84", X"13",
     X"24", X"d6", X"10", X"08", X"68", X"68", X"20", X"65",
     X"d6", X"4c", X"d2", X"d7", X"e8", X"bd", X"00", X"02",
     X"24", X"13", X"70", X"04", X"c9", X"20", X"f0", X"f4",
     X"85", X"0e", X"c9", X"22", X"f0", X"74", X"70", X"4d",
     X"c9", X"3f", X"d0", X"04", X"a9", X"ba", X"d0", X"45",
     X"c9", X"30", X"90", X"04", X"c9", X"3c", X"90", X"3d",
     X"84", X"ad", X"a9", X"d0", X"85", X"9d", X"a9", X"cf",
     X"85", X"9e", X"a0", X"00", X"84", X"0f", X"88", X"86",
     X"b8", X"ca", X"c8", X"d0", X"02", X"e6", X"9e", X"e8",
     X"bd", X"00", X"02", X"c9", X"20", X"f0", X"f8", X"38",
     X"f1", X"9d", X"f0", X"ee", X"c9", X"80", X"d0", X"41",
     X"05", X"0f", X"c9", X"c5", X"d0", X"0d", X"bd", X"01",
     X"02", X"c9", X"4e", X"f0", X"34", X"c9", X"4f", X"f0",
     X"30", X"a9", X"c5", X"a4", X"ad", X"e8", X"c8", X"99",
     X"fb", X"01", X"b9", X"fb", X"01", X"f0", X"39", X"38",
     X"e9", X"3a", X"f0", X"04", X"c9", X"49", X"d0", X"02",
     X"85", X"13", X"38", X"e9", X"78", X"d0", X"86", X"85",
     X"0e", X"bd", X"00", X"02", X"f0", X"df", X"c5", X"0e",
     X"f0", X"db", X"c8", X"99", X"fb", X"01", X"e8", X"d0",
     X"f0", X"a6", X"b8", X"e6", X"0f", X"b1", X"9d", X"c8",
     X"d0", X"02", X"e6", X"9e", X"0a", X"90", X"f6", X"b1",
     X"9d", X"d0", X"9d", X"bd", X"00", X"02", X"10", X"bb",
     X"99", X"fd", X"01", X"c6", X"b9", X"a9", X"ff", X"85",
     X"b8", X"60", X"a5", X"67", X"a6", X"68", X"a0", X"01",
     X"85", X"9b", X"86", X"9c", X"b1", X"9b", X"f0", X"1f",
     X"c8", X"c8", X"a5", X"51", X"d1", X"9b", X"90", X"18",
     X"f0", X"03", X"88", X"d0", X"09", X"a5", X"50", X"88",
     X"d1", X"9b", X"90", X"0c", X"f0", X"0a", X"88", X"b1",
     X"9b", X"aa", X"88", X"b1", X"9b", X"b0", X"d7", X"18",
     X"60", X"d0", X"fd", X"a9", X"00", X"85", X"d6", X"a8",
     X"91", X"67", X"c8", X"91", X"67", X"a5", X"67", X"69",
     X"02", X"85", X"69", X"85", X"af", X"a5", X"68", X"69",
     X"00", X"85", X"6a", X"85", X"b0", X"20", X"97", X"d6",
     X"a9", X"00", X"d0", X"2a", X"a5", X"73", X"a4", X"74",
     X"85", X"6f", X"84", X"70", X"a5", X"69", X"a4", X"6a",
     X"85", X"6b", X"84", X"6c", X"85", X"6d", X"84", X"6e",
     X"20", X"49", X"d8", X"a2", X"55", X"86", X"52", X"68",
     X"a8", X"68", X"a2", X"f8", X"9a", X"48", X"98", X"48",
     X"a9", X"00", X"85", X"7a", X"85", X"14", X"60", X"18",
     X"a5", X"67", X"69", X"ff", X"85", X"b8", X"a5", X"68",
     X"69", X"ff", X"85", X"b9", X"60", X"90", X"0a", X"f0",
     X"08", X"c9", X"c9", X"f0", X"04", X"c9", X"2c", X"d0",
     X"e5", X"20", X"0c", X"da", X"20", X"1a", X"d6", X"20",
     X"b7", X"00", X"f0", X"10", X"c9", X"c9", X"f0", X"04",
     X"c9", X"2c", X"d0", X"84", X"20", X"b1", X"00", X"20",
     X"0c", X"da", X"d0", X"ca", X"68", X"68", X"a5", X"50",
     X"05", X"51", X"d0", X"06", X"a9", X"ff", X"85", X"50",
     X"85", X"51", X"a0", X"01", X"b1", X"9b", X"f0", X"44",
     X"20", X"58", X"d8", X"20", X"fb", X"da", X"c8", X"b1",
     X"9b", X"aa", X"c8", X"b1", X"9b", X"c5", X"51", X"d0",
     X"04", X"e4", X"50", X"f0", X"02", X"b0", X"2d", X"84",
     X"85", X"20", X"24", X"ed", X"a9", X"20", X"a4", X"85",
     X"29", X"7f", X"20", X"5c", X"db", X"a5", X"24", X"c9",
     X"21", X"90", X"07", X"20", X"fb", X"da", X"a9", X"05",
     X"85", X"24", X"c8", X"b1", X"9b", X"d0", X"1d", X"a8",
     X"b1", X"9b", X"aa", X"c8", X"b1", X"9b", X"86", X"9b",
     X"85", X"9c", X"d0", X"b6", X"a9", X"0d", X"20", X"5c",
     X"db", X"4c", X"d2", X"d7", X"c8", X"d0", X"02", X"e6",
     X"9e", X"b1", X"9d", X"60", X"10", X"cc", X"38", X"e9",
     X"7f", X"aa", X"84", X"85", X"a0", X"d0", X"84", X"9d",
     X"a0", X"cf", X"84", X"9e", X"a0", X"ff", X"ca", X"f0",
     X"07", X"20", X"2c", X"d7", X"10", X"fb", X"30", X"f6",
     X"a9", X"20", X"20", X"5c", X"db", X"20", X"2c", X"d7",
     X"30", X"05", X"20", X"5c", X"db", X"d0", X"f6", X"20",
     X"5c", X"db", X"a9", X"20", X"d0", X"98", X"a9", X"80",
     X"85", X"14", X"20", X"46", X"da", X"20", X"65", X"d3",
     X"d0", X"05", X"8a", X"69", X"0f", X"aa", X"9a", X"68",
     X"68", X"a9", X"09", X"20", X"d6", X"d3", X"20", X"a3",
     X"d9", X"18", X"98", X"65", X"b8", X"48", X"a5", X"b9",
     X"69", X"00", X"48", X"a5", X"76", X"48", X"a5", X"75",
     X"48", X"a9", X"c1", X"20", X"c0", X"de", X"20", X"6a",
     X"dd", X"20", X"67", X"dd", X"a5", X"a2", X"09", X"7f",
     X"25", X"9e", X"85", X"9e", X"a9", X"af", X"a0", X"d7",
     X"85", X"5e", X"84", X"5f", X"4c", X"20", X"de", X"a9",
     X"13", X"a0", X"e9", X"20", X"f9", X"ea", X"20", X"b7",
     X"00", X"c9", X"c7", X"d0", X"06", X"20", X"b1", X"00",
     X"20", X"67", X"dd", X"20", X"82", X"eb", X"20", X"15",
     X"de", X"a5", X"86", X"48", X"a5", X"85", X"48", X"a9",
     X"81", X"48", X"ba", X"86", X"f8", X"20", X"58", X"d8",
     X"a5", X"b8", X"a4", X"b9", X"a6", X"76", X"e8", X"f0",
     X"04", X"85", X"79", X"84", X"7a", X"a0", X"00", X"b1",
     X"b8", X"d0", X"57", X"a0", X"02", X"b1", X"b8", X"18",
     X"f0", X"34", X"c8", X"b1", X"b8", X"85", X"75", X"c8",
     X"b1", X"b8", X"85", X"76", X"98", X"65", X"b8", X"85",
     X"b8", X"90", X"02", X"e6", X"b9", X"24", X"f2", X"10",
     X"14", X"a6", X"76", X"e8", X"f0", X"0f", X"a9", X"23",
     X"20", X"5c", X"db", X"a6", X"75", X"a5", X"76", X"20",
     X"24", X"ed", X"20", X"57", X"db", X"20", X"b1", X"00",
     X"20", X"28", X"d8", X"4c", X"d2", X"d7", X"f0", X"62",
     X"f0", X"2d", X"e9", X"80", X"90", X"11", X"c9", X"40",
     X"b0", X"14", X"0a", X"a8", X"b9", X"01", X"d0", X"48",
     X"b9", X"00", X"d0", X"48", X"4c", X"b1", X"00", X"4c",
     X"46", X"da", X"c9", X"3a", X"f0", X"bf", X"4c", X"c9",
     X"de", X"38", X"a5", X"67", X"e9", X"01", X"a4", X"68",
     X"b0", X"01", X"88", X"85", X"7d", X"84", X"7e", X"60",
     X"ad", X"00", X"c0", X"c9", X"83", X"f0", X"01", X"60",
     X"20", X"53", X"d5", X"a2", X"ff", X"24", X"d8", X"10",
     X"03", X"4c", X"e9", X"f2", X"c9", X"03", X"b0", X"01",
     X"18", X"d0", X"3c", X"a5", X"b8", X"a4", X"b9", X"a6",
     X"76", X"e8", X"f0", X"0c", X"85", X"79", X"84", X"7a",
     X"a5", X"75", X"a4", X"76", X"85", X"77", X"84", X"78",
     X"68", X"68", X"a9", X"5d", X"a0", X"d3", X"90", X"03",
     X"4c", X"31", X"d4", X"4c", X"3c", X"d4", X"d0", X"17",
     X"a2", X"d2", X"a4", X"7a", X"d0", X"03", X"4c", X"12",
     X"d4", X"a5", X"79", X"85", X"b8", X"84", X"b9", X"a5",
     X"77", X"a4", X"78", X"85", X"75", X"84", X"76", X"60",
     X"38", X"a5", X"af", X"e5", X"67", X"85", X"50", X"a5",
     X"b0", X"e5", X"68", X"85", X"51", X"20", X"f0", X"d8",
     X"20", X"cd", X"fe", X"20", X"01", X"d9", X"4c", X"cd",
     X"fe", X"20", X"f0", X"d8", X"20", X"fd", X"fe", X"18",
     X"a5", X"67", X"65", X"50", X"85", X"69", X"a5", X"68",
     X"65", X"51", X"85", X"6a", X"a5", X"52", X"85", X"d6",
     X"20", X"01", X"d9", X"20", X"fd", X"fe", X"24", X"d6",
     X"10", X"03", X"4c", X"65", X"d6", X"4c", X"f2", X"d4",
     X"a9", X"50", X"a0", X"00", X"85", X"3c", X"84", X"3d",
     X"a9", X"52", X"85", X"3e", X"84", X"3f", X"84", X"d6",
     X"60", X"a5", X"67", X"a4", X"68", X"85", X"3c", X"84",
     X"3d", X"a5", X"69", X"a4", X"6a", X"85", X"3e", X"84",
     X"3f", X"60", X"08", X"c6", X"76", X"28", X"d0", X"03",
     X"4c", X"65", X"d6", X"20", X"6c", X"d6", X"4c", X"35",
     X"d9", X"a9", X"03", X"20", X"d6", X"d3", X"a5", X"b9",
     X"48", X"a5", X"b8", X"48", X"a5", X"76", X"48", X"a5",
     X"75", X"48", X"a9", X"b0", X"48", X"20", X"b7", X"00",
     X"20", X"3e", X"d9", X"4c", X"d2", X"d7", X"20", X"0c",
     X"da", X"20", X"a6", X"d9", X"a5", X"76", X"c5", X"51",
     X"b0", X"0b", X"98", X"38", X"65", X"b8", X"a6", X"b9",
     X"90", X"07", X"e8", X"b0", X"04", X"a5", X"67", X"a6",
     X"68", X"20", X"1e", X"d6", X"90", X"1e", X"a5", X"9b",
     X"e9", X"01", X"85", X"b8", X"a5", X"9c", X"e9", X"00",
     X"85", X"b9", X"60", X"d0", X"fd", X"a9", X"ff", X"85",
     X"85", X"20", X"65", X"d3", X"9a", X"c9", X"b0", X"f0",
     X"0b", X"a2", X"16", X"2c", X"a2", X"5a", X"4c", X"12",
     X"d4", X"4c", X"c9", X"de", X"68", X"68", X"c0", X"42",
     X"f0", X"3b", X"85", X"75", X"68", X"85", X"76", X"68",
     X"85", X"b8", X"68", X"85", X"b9", X"20", X"a3", X"d9",
     X"98", X"18", X"65", X"b8", X"85", X"b8", X"90", X"02",
     X"e6", X"b9", X"60", X"a2", X"3a", X"2c", X"a2", X"00",
     X"86", X"0d", X"a0", X"00", X"84", X"0e", X"a5", X"0e",
     X"a6", X"0d", X"85", X"0d", X"86", X"0e", X"b1", X"b8",
     X"f0", X"e8", X"c5", X"0e", X"f0", X"e4", X"c8", X"c9",
     X"22", X"d0", X"f3", X"f0", X"e9", X"68", X"68", X"68",
     X"60", X"20", X"7b", X"dd", X"20", X"b7", X"00", X"c9",
     X"ab", X"f0", X"05", X"a9", X"c4", X"20", X"c0", X"de",
     X"a5", X"9d", X"d0", X"05", X"20", X"a6", X"d9", X"f0",
     X"b7", X"20", X"b7", X"00", X"b0", X"03", X"4c", X"3e",
     X"d9", X"4c", X"28", X"d8", X"20", X"f8", X"e6", X"48",
     X"c9", X"b0", X"f0", X"04", X"c9", X"ab", X"d0", X"89",
     X"c6", X"a1", X"d0", X"04", X"68", X"4c", X"2a", X"d8",
     X"20", X"b1", X"00", X"20", X"0c", X"da", X"c9", X"2c",
     X"f0", X"ee", X"68", X"60", X"a2", X"00", X"86", X"50",
     X"86", X"51", X"b0", X"f7", X"e9", X"2f", X"85", X"0d",
     X"a5", X"51", X"85", X"5e", X"c9", X"19", X"b0", X"d4",
     X"a5", X"50", X"0a", X"26", X"5e", X"0a", X"26", X"5e",
     X"65", X"50", X"85", X"50", X"a5", X"5e", X"65", X"51",
     X"85", X"51", X"06", X"50", X"26", X"51", X"a5", X"50",
     X"65", X"0d", X"85", X"50", X"90", X"02", X"e6", X"51",
     X"20", X"b1", X"00", X"4c", X"12", X"da", X"20", X"e3",
     X"df", X"85", X"85", X"84", X"86", X"a9", X"d0", X"20",
     X"c0", X"de", X"a5", X"12", X"48", X"a5", X"11", X"48",
     X"20", X"7b", X"dd", X"68", X"2a", X"20", X"6d", X"dd",
     X"d0", X"18", X"68", X"10", X"12", X"20", X"72", X"eb",
     X"20", X"0c", X"e1", X"a0", X"00", X"a5", X"a0", X"91",
     X"85", X"c8", X"a5", X"a1", X"91", X"85", X"60", X"4c",
     X"27", X"eb", X"68", X"a0", X"02", X"b1", X"a0", X"c5",
     X"70", X"90", X"17", X"d0", X"07", X"88", X"b1", X"a0",
     X"c5", X"6f", X"90", X"0e", X"a4", X"a1", X"c4", X"6a",
     X"90", X"08", X"d0", X"0d", X"a5", X"a0", X"c5", X"69",
     X"b0", X"07", X"a5", X"a0", X"a4", X"a1", X"4c", X"b7",
     X"da", X"a0", X"00", X"b1", X"a0", X"20", X"d5", X"e3",
     X"a5", X"8c", X"a4", X"8d", X"85", X"ab", X"84", X"ac",
     X"20", X"d4", X"e5", X"a9", X"9d", X"a0", X"00", X"85",
     X"8c", X"84", X"8d", X"20", X"35", X"e6", X"a0", X"00",
     X"b1", X"8c", X"91", X"85", X"c8", X"b1", X"8c", X"91",
     X"85", X"c8", X"b1", X"8c", X"91", X"85", X"60", X"20",
     X"3d", X"db", X"20", X"b7", X"00", X"f0", X"24", X"f0",
     X"29", X"c9", X"c0", X"f0", X"39", X"c9", X"c3", X"18",
     X"f0", X"34", X"c9", X"2c", X"18", X"f0", X"1c", X"c9",
     X"3b", X"f0", X"44", X"20", X"7b", X"dd", X"24", X"11",
     X"30", X"dd", X"20", X"34", X"ed", X"20", X"e7", X"e3",
     X"4c", X"cf", X"da", X"a9", X"0d", X"20", X"5c", X"db",
     X"49", X"ff", X"60", X"a5", X"24", X"c9", X"18", X"90",
     X"05", X"20", X"fb", X"da", X"d0", X"21", X"69", X"10",
     X"29", X"f0", X"85", X"24", X"90", X"19", X"08", X"20",
     X"f5", X"e6", X"c9", X"29", X"f0", X"03", X"4c", X"c9",
     X"de", X"28", X"90", X"07", X"ca", X"8a", X"e5", X"24",
     X"90", X"05", X"aa", X"e8", X"ca", X"d0", X"06", X"20",
     X"b1", X"00", X"4c", X"d7", X"da", X"20", X"57", X"db",
     X"d0", X"f2", X"20", X"e7", X"e3", X"20", X"00", X"e6",
     X"aa", X"a0", X"00", X"e8", X"ca", X"f0", X"bb", X"b1",
     X"5e", X"20", X"5c", X"db", X"c8", X"c9", X"0d", X"d0",
     X"f3", X"20", X"00", X"db", X"4c", X"44", X"db", X"a9",
     X"20", X"2c", X"a9", X"3f", X"09", X"80", X"c9", X"a0",
     X"90", X"02", X"05", X"f3", X"20", X"ed", X"fd", X"29",
     X"7f", X"48", X"a5", X"f1", X"20", X"a8", X"fc", X"68",
     X"60", X"a5", X"15", X"f0", X"12", X"30", X"04", X"a0",
     X"ff", X"d0", X"04", X"a5", X"7b", X"a4", X"7c", X"85",
     X"75", X"84", X"76", X"4c", X"c9", X"de", X"68", X"24",
     X"d8", X"10", X"05", X"a2", X"fe", X"4c", X"e9", X"f2",
     X"a9", X"ef", X"a0", X"dc", X"20", X"3a", X"db", X"a5",
     X"79", X"a4", X"7a", X"85", X"b8", X"84", X"b9", X"60",
     X"20", X"06", X"e3", X"a2", X"01", X"a0", X"02", X"a9",
     X"00", X"8d", X"01", X"02", X"a9", X"40", X"20", X"eb",
     X"db", X"60", X"c9", X"22", X"d0", X"0e", X"20", X"81",
     X"de", X"a9", X"3b", X"20", X"c0", X"de", X"20", X"3d",
     X"db", X"4c", X"c7", X"db", X"20", X"5a", X"db", X"20",
     X"06", X"e3", X"a9", X"2c", X"8d", X"ff", X"01", X"20",
     X"2c", X"d5", X"ad", X"00", X"02", X"c9", X"03", X"d0",
     X"10", X"4c", X"63", X"d8", X"20", X"5a", X"db", X"4c",
     X"2c", X"d5", X"a6", X"7d", X"a4", X"7e", X"a9", X"98",
     X"2c", X"a9", X"00", X"85", X"15", X"86", X"7f", X"84",
     X"80", X"20", X"e3", X"df", X"85", X"85", X"84", X"86",
     X"a5", X"b8", X"a4", X"b9", X"85", X"87", X"84", X"88",
     X"a6", X"7f", X"a4", X"80", X"86", X"b8", X"84", X"b9",
     X"20", X"b7", X"00", X"d0", X"1e", X"24", X"15", X"50",
     X"0e", X"20", X"0c", X"fd", X"29", X"7f", X"8d", X"00",
     X"02", X"a2", X"ff", X"a0", X"01", X"d0", X"08", X"30",
     X"7f", X"20", X"5a", X"db", X"20", X"dc", X"db", X"86",
     X"b8", X"84", X"b9", X"20", X"b1", X"00", X"24", X"11",
     X"10", X"31", X"24", X"15", X"50", X"09", X"e8", X"86",
     X"b8", X"a9", X"00", X"85", X"0d", X"f0", X"0c", X"85",
     X"0d", X"c9", X"22", X"f0", X"07", X"a9", X"3a", X"85",
     X"0d", X"a9", X"2c", X"18", X"85", X"0e", X"a5", X"b8",
     X"a4", X"b9", X"69", X"00", X"90", X"01", X"c8", X"20",
     X"ed", X"e3", X"20", X"3d", X"e7", X"20", X"7b", X"da",
     X"4c", X"72", X"dc", X"48", X"ad", X"00", X"02", X"f0",
     X"30", X"68", X"20", X"4a", X"ec", X"a5", X"12", X"20",
     X"63", X"da", X"20", X"b7", X"00", X"f0", X"07", X"c9",
     X"2c", X"f0", X"03", X"4c", X"71", X"db", X"a5", X"b8",
     X"a4", X"b9", X"85", X"7f", X"84", X"80", X"a5", X"87",
     X"a4", X"88", X"85", X"b8", X"84", X"b9", X"20", X"b7",
     X"00", X"f0", X"33", X"20", X"be", X"de", X"4c", X"f1",
     X"db", X"a5", X"15", X"d0", X"cc", X"4c", X"86", X"db",
     X"20", X"a3", X"d9", X"c8", X"aa", X"d0", X"12", X"a2",
     X"2a", X"c8", X"b1", X"b8", X"f0", X"5f", X"c8", X"b1",
     X"b8", X"85", X"7b", X"c8", X"b1", X"b8", X"c8", X"85",
     X"7c", X"b1", X"b8", X"aa", X"20", X"98", X"d9", X"e0",
     X"83", X"d0", X"dd", X"4c", X"2b", X"dc", X"a5", X"7f",
     X"a4", X"80", X"a6", X"15", X"10", X"03", X"4c", X"53",
     X"d8", X"a0", X"00", X"b1", X"7f", X"f0", X"07", X"a9",
     X"df", X"a0", X"dc", X"4c", X"3a", X"db", X"60", X"3f",
     X"45", X"58", X"54", X"52", X"41", X"20", X"49", X"47",
     X"4e", X"4f", X"52", X"45", X"44", X"0d", X"00", X"3f",
     X"52", X"45", X"45", X"4e", X"54", X"45", X"52", X"0d",
     X"00", X"d0", X"04", X"a0", X"00", X"f0", X"03", X"20",
     X"e3", X"df", X"85", X"85", X"84", X"86", X"20", X"65",
     X"d3", X"f0", X"04", X"a2", X"00", X"f0", X"69", X"9a",
     X"e8", X"e8", X"e8", X"e8", X"8a", X"e8", X"e8", X"e8",
     X"e8", X"e8", X"e8", X"86", X"60", X"a0", X"01", X"20",
     X"f9", X"ea", X"ba", X"bd", X"09", X"01", X"85", X"a2",
     X"a5", X"85", X"a4", X"86", X"20", X"be", X"e7", X"20",
     X"27", X"eb", X"a0", X"01", X"20", X"b4", X"eb", X"ba",
     X"38", X"fd", X"09", X"01", X"f0", X"17", X"bd", X"0f",
     X"01", X"85", X"75", X"bd", X"10", X"01", X"85", X"76",
     X"bd", X"12", X"01", X"85", X"b8", X"bd", X"11", X"01",
     X"85", X"b9", X"4c", X"d2", X"d7", X"8a", X"69", X"11",
     X"aa", X"9a", X"20", X"b7", X"00", X"c9", X"2c", X"d0",
     X"f1", X"20", X"b1", X"00", X"20", X"ff", X"dc", X"20",
     X"7b", X"dd", X"18", X"24", X"38", X"24", X"11", X"30",
     X"03", X"b0", X"03", X"60", X"b0", X"fd", X"a2", X"a3",
     X"4c", X"12", X"d4", X"a6", X"b8", X"d0", X"02", X"c6",
     X"b9", X"c6", X"b8", X"a2", X"00", X"24", X"48", X"8a",
     X"48", X"a9", X"01", X"20", X"d6", X"d3", X"20", X"60",
     X"de", X"a9", X"00", X"85", X"89", X"20", X"b7", X"00",
     X"38", X"e9", X"cf", X"90", X"17", X"c9", X"03", X"b0",
     X"13", X"c9", X"01", X"2a", X"49", X"01", X"45", X"89",
     X"c5", X"89", X"90", X"61", X"85", X"89", X"20", X"b1",
     X"00", X"4c", X"98", X"dd", X"a6", X"89", X"d0", X"2c",
     X"b0", X"7b", X"69", X"07", X"90", X"77", X"65", X"11",
     X"d0", X"03", X"4c", X"97", X"e5", X"69", X"ff", X"85",
     X"5e", X"0a", X"65", X"5e", X"a8", X"68", X"d9", X"b2",
     X"d0", X"b0", X"67", X"20", X"6a", X"dd", X"48", X"20",
     X"fd", X"dd", X"68", X"a4", X"87", X"10", X"17", X"aa",
     X"f0", X"56", X"d0", X"5f", X"46", X"11", X"8a", X"2a",
     X"a6", X"b8", X"d0", X"02", X"c6", X"b9", X"c6", X"b8",
     X"a0", X"1b", X"85", X"89", X"d0", X"d7", X"d9", X"b2",
     X"d0", X"b0", X"48", X"90", X"d9", X"b9", X"b4", X"d0",
     X"48", X"b9", X"b3", X"d0", X"48", X"20", X"10", X"de",
     X"a5", X"89", X"4c", X"86", X"dd", X"4c", X"c9", X"de",
     X"a5", X"a2", X"be", X"b2", X"d0", X"a8", X"68", X"85",
     X"5e", X"e6", X"5e", X"68", X"85", X"5f", X"98", X"48",
     X"20", X"72", X"eb", X"a5", X"a1", X"48", X"a5", X"a0",
     X"48", X"a5", X"9f", X"48", X"a5", X"9e", X"48", X"a5",
     X"9d", X"48", X"6c", X"5e", X"00", X"a0", X"ff", X"68",
     X"f0", X"23", X"c9", X"64", X"f0", X"03", X"20", X"6a",
     X"dd", X"84", X"87", X"68", X"4a", X"85", X"16", X"68",
     X"85", X"a5", X"68", X"85", X"a6", X"68", X"85", X"a7",
     X"68", X"85", X"a8", X"68", X"85", X"a9", X"68", X"85",
     X"aa", X"45", X"a2", X"85", X"ab", X"a5", X"9d", X"60",
     X"a9", X"00", X"85", X"11", X"20", X"b1", X"00", X"b0",
     X"03", X"4c", X"4a", X"ec", X"20", X"7d", X"e0", X"b0",
     X"64", X"c9", X"2e", X"f0", X"f4", X"c9", X"c9", X"f0",
     X"55", X"c9", X"c8", X"f0", X"e7", X"c9", X"22", X"d0",
     X"0f", X"a5", X"b8", X"a4", X"b9", X"69", X"00", X"90",
     X"01", X"c8", X"20", X"e7", X"e3", X"4c", X"3d", X"e7",
     X"c9", X"c6", X"d0", X"10", X"a0", X"18", X"d0", X"38",
     X"a5", X"9d", X"d0", X"03", X"a0", X"01", X"2c", X"a0",
     X"00", X"4c", X"01", X"e3", X"c9", X"c2", X"d0", X"03",
     X"4c", X"54", X"e3", X"c9", X"d2", X"90", X"03", X"4c",
     X"0c", X"df", X"20", X"bb", X"de", X"20", X"7b", X"dd",
     X"a9", X"29", X"2c", X"a9", X"28", X"2c", X"a9", X"2c",
     X"a0", X"00", X"d1", X"b8", X"d0", X"03", X"4c", X"b1",
     X"00", X"a2", X"10", X"4c", X"12", X"d4", X"a0", X"15",
     X"68", X"68", X"4c", X"d7", X"dd", X"20", X"e3", X"df",
     X"85", X"a0", X"84", X"a1", X"a6", X"11", X"f0", X"05",
     X"a2", X"00", X"86", X"ac", X"60", X"a6", X"12", X"10",
     X"0d", X"a0", X"00", X"b1", X"a0", X"aa", X"c8", X"b1",
     X"a0", X"a8", X"8a", X"4c", X"f2", X"e2", X"4c", X"f9",
     X"ea", X"20", X"b1", X"00", X"20", X"ec", X"f1", X"8a",
     X"a4", X"f0", X"20", X"71", X"f8", X"a8", X"20", X"01",
     X"e3", X"4c", X"b8", X"de", X"c9", X"d7", X"f0", X"e9",
     X"0a", X"48", X"aa", X"20", X"b1", X"00", X"e0", X"cf",
     X"90", X"20", X"20", X"bb", X"de", X"20", X"7b", X"dd",
     X"20", X"be", X"de", X"20", X"6c", X"dd", X"68", X"aa",
     X"a5", X"a1", X"48", X"a5", X"a0", X"48", X"8a", X"48",
     X"20", X"f8", X"e6", X"68", X"a8", X"8a", X"48", X"4c",
     X"3f", X"df", X"20", X"b2", X"de", X"68", X"a8", X"b9",
     X"dc", X"cf", X"85", X"91", X"b9", X"dd", X"cf", X"85",
     X"92", X"20", X"90", X"00", X"4c", X"6a", X"dd", X"a5",
     X"a5", X"05", X"9d", X"d0", X"0b", X"a5", X"a5", X"f0",
     X"04", X"a5", X"9d", X"d0", X"03", X"a0", X"00", X"2c",
     X"a0", X"01", X"4c", X"01", X"e3", X"20", X"6d", X"dd",
     X"b0", X"13", X"a5", X"aa", X"09", X"7f", X"25", X"a6",
     X"85", X"a6", X"a9", X"a5", X"a0", X"00", X"20", X"b2",
     X"eb", X"aa", X"4c", X"b0", X"df", X"a9", X"00", X"85",
     X"11", X"c6", X"89", X"20", X"00", X"e6", X"85", X"9d",
     X"86", X"9e", X"84", X"9f", X"a5", X"a8", X"a4", X"a9",
     X"20", X"04", X"e6", X"86", X"a8", X"84", X"a9", X"aa",
     X"38", X"e5", X"9d", X"f0", X"08", X"a9", X"01", X"90",
     X"04", X"a6", X"9d", X"a9", X"ff", X"85", X"a2", X"a0",
     X"ff", X"e8", X"c8", X"ca", X"d0", X"07", X"a6", X"a2",
     X"30", X"0f", X"18", X"90", X"0c", X"b1", X"a8", X"d1",
     X"9e", X"f0", X"ef", X"a2", X"ff", X"b0", X"02", X"a2",
     X"01", X"e8", X"8a", X"2a", X"25", X"16", X"f0", X"02",
     X"a9", X"01", X"4c", X"93", X"eb", X"20", X"fb", X"e6",
     X"20", X"1e", X"fb", X"4c", X"01", X"e3", X"20", X"be",
     X"de", X"aa", X"20", X"e8", X"df", X"20", X"b7", X"00",
     X"d0", X"f4", X"60", X"a2", X"00", X"20", X"b7", X"00",
     X"86", X"10", X"85", X"81", X"20", X"b7", X"00", X"20",
     X"7d", X"e0", X"b0", X"03", X"4c", X"c9", X"de", X"a2",
     X"00", X"86", X"11", X"86", X"12", X"4c", X"07", X"e0",
     X"4c", X"28", X"f1", X"4c", X"3c", X"d4", X"00", X"20",
     X"b1", X"00", X"90", X"05", X"20", X"7d", X"e0", X"90",
     X"0b", X"aa", X"20", X"b1", X"00", X"90", X"fb", X"20",
     X"7d", X"e0", X"b0", X"f6", X"c9", X"24", X"d0", X"06",
     X"a9", X"ff", X"85", X"11", X"d0", X"10", X"c9", X"25",
     X"d0", X"13", X"a5", X"14", X"30", X"c6", X"a9", X"80",
     X"85", X"12", X"05", X"81", X"85", X"81", X"8a", X"09",
     X"80", X"aa", X"20", X"b1", X"00", X"86", X"82", X"38",
     X"05", X"14", X"e9", X"28", X"d0", X"03", X"4c", X"1e",
     X"e1", X"24", X"14", X"30", X"02", X"70", X"f7", X"a9",
     X"00", X"85", X"14", X"a5", X"69", X"a6", X"6a", X"a0",
     X"00", X"86", X"9c", X"85", X"9b", X"e4", X"6c", X"d0",
     X"04", X"c5", X"6b", X"f0", X"22", X"a5", X"81", X"d1",
     X"9b", X"d0", X"08", X"a5", X"82", X"c8", X"d1", X"9b",
     X"f0", X"6c", X"88", X"18", X"a5", X"9b", X"69", X"07",
     X"90", X"e1", X"e8", X"d0", X"dc", X"c9", X"41", X"90",
     X"05", X"e9", X"5b", X"38", X"e9", X"a5", X"60", X"68",
     X"48", X"c9", X"d7", X"d0", X"0f", X"ba", X"bd", X"02",
     X"01", X"c9", X"de", X"d0", X"07", X"a9", X"9a", X"a0",
     X"e0", X"60", X"00", X"00", X"a5", X"6b", X"a4", X"6c",
     X"85", X"9b", X"84", X"9c", X"a5", X"6d", X"a4", X"6e",
     X"85", X"96", X"84", X"97", X"18", X"69", X"07", X"90",
     X"01", X"c8", X"85", X"94", X"84", X"95", X"20", X"93",
     X"d3", X"a5", X"94", X"a4", X"95", X"c8", X"85", X"6b",
     X"84", X"6c", X"a0", X"00", X"a5", X"81", X"91", X"9b",
     X"c8", X"a5", X"82", X"91", X"9b", X"a9", X"00", X"c8",
     X"91", X"9b", X"c8", X"91", X"9b", X"c8", X"91", X"9b",
     X"c8", X"91", X"9b", X"c8", X"91", X"9b", X"a5", X"9b",
     X"18", X"69", X"02", X"a4", X"9c", X"90", X"01", X"c8",
     X"85", X"83", X"84", X"84", X"60", X"a5", X"0f", X"0a",
     X"69", X"05", X"65", X"9b", X"a4", X"9c", X"90", X"01",
     X"c8", X"85", X"94", X"84", X"95", X"60", X"90", X"80",
     X"00", X"00", X"20", X"b1", X"00", X"20", X"67", X"dd",
     X"a5", X"a2", X"30", X"0d", X"a5", X"9d", X"c9", X"90",
     X"90", X"09", X"a9", X"fe", X"a0", X"e0", X"20", X"b2",
     X"eb", X"d0", X"7e", X"4c", X"f2", X"eb", X"a5", X"14",
     X"d0", X"47", X"a5", X"10", X"05", X"12", X"48", X"a5",
     X"11", X"48", X"a0", X"00", X"98", X"48", X"a5", X"82",
     X"48", X"a5", X"81", X"48", X"20", X"02", X"e1", X"68",
     X"85", X"81", X"68", X"85", X"82", X"68", X"a8", X"ba",
     X"bd", X"02", X"01", X"48", X"bd", X"01", X"01", X"48",
     X"a5", X"a0", X"9d", X"02", X"01", X"a5", X"a1", X"9d",
     X"01", X"01", X"c8", X"20", X"b7", X"00", X"c9", X"2c",
     X"f0", X"d2", X"84", X"0f", X"20", X"b8", X"de", X"68",
     X"85", X"11", X"68", X"85", X"12", X"29", X"7f", X"85",
     X"10", X"a6", X"6b", X"a5", X"6c", X"86", X"9b", X"85",
     X"9c", X"c5", X"6e", X"d0", X"04", X"e4", X"6d", X"f0",
     X"3f", X"a0", X"00", X"b1", X"9b", X"c8", X"c5", X"81",
     X"d0", X"06", X"a5", X"82", X"d1", X"9b", X"f0", X"16",
     X"c8", X"b1", X"9b", X"18", X"65", X"9b", X"aa", X"c8",
     X"b1", X"9b", X"65", X"9c", X"90", X"d7", X"a2", X"6b",
     X"2c", X"a2", X"35", X"4c", X"12", X"d4", X"a2", X"78",
     X"a5", X"10", X"d0", X"f7", X"a5", X"14", X"f0", X"02",
     X"38", X"60", X"20", X"ed", X"e0", X"a5", X"0f", X"a0",
     X"04", X"d1", X"9b", X"d0", X"e1", X"4c", X"4b", X"e2",
     X"a5", X"14", X"f0", X"05", X"a2", X"2a", X"4c", X"12",
     X"d4", X"20", X"ed", X"e0", X"20", X"e3", X"d3", X"a9",
     X"00", X"a8", X"85", X"ae", X"a2", X"05", X"a5", X"81",
     X"91", X"9b", X"10", X"01", X"ca", X"c8", X"a5", X"82",
     X"91", X"9b", X"10", X"02", X"ca", X"ca", X"86", X"ad",
     X"a5", X"0f", X"c8", X"c8", X"c8", X"91", X"9b", X"a2",
     X"0b", X"a9", X"00", X"24", X"10", X"50", X"08", X"68",
     X"18", X"69", X"01", X"aa", X"68", X"69", X"00", X"c8",
     X"91", X"9b", X"c8", X"8a", X"91", X"9b", X"20", X"ad",
     X"e2", X"86", X"ad", X"85", X"ae", X"a4", X"5e", X"c6",
     X"0f", X"d0", X"dc", X"65", X"95", X"b0", X"5d", X"85",
     X"95", X"a8", X"8a", X"65", X"94", X"90", X"03", X"c8",
     X"f0", X"52", X"20", X"e3", X"d3", X"85", X"6d", X"84",
     X"6e", X"a9", X"00", X"e6", X"ae", X"a4", X"ad", X"f0",
     X"05", X"88", X"91", X"94", X"d0", X"fb", X"c6", X"95",
     X"c6", X"ae", X"d0", X"f5", X"e6", X"95", X"38", X"a5",
     X"6d", X"e5", X"9b", X"a0", X"02", X"91", X"9b", X"a5",
     X"6e", X"c8", X"e5", X"9c", X"91", X"9b", X"a5", X"10",
     X"d0", X"62", X"c8", X"b1", X"9b", X"85", X"0f", X"a9",
     X"00", X"85", X"ad", X"85", X"ae", X"c8", X"68", X"aa",
     X"85", X"a0", X"68", X"85", X"a1", X"d1", X"9b", X"90",
     X"0e", X"d0", X"06", X"c8", X"8a", X"d1", X"9b", X"90",
     X"07", X"4c", X"96", X"e1", X"4c", X"10", X"d4", X"c8",
     X"a5", X"ae", X"05", X"ad", X"18", X"f0", X"0a", X"20",
     X"ad", X"e2", X"8a", X"65", X"a0", X"aa", X"98", X"a4",
     X"5e", X"65", X"a1", X"86", X"ad", X"c6", X"0f", X"d0",
     X"ca", X"85", X"ae", X"a2", X"05", X"a5", X"81", X"10",
     X"01", X"ca", X"a5", X"82", X"10", X"02", X"ca", X"ca",
     X"86", X"64", X"a9", X"00", X"20", X"b6", X"e2", X"8a",
     X"65", X"94", X"85", X"83", X"98", X"65", X"95", X"85",
     X"84", X"a8", X"a5", X"83", X"60", X"84", X"5e", X"b1",
     X"9b", X"85", X"64", X"88", X"b1", X"9b", X"85", X"65",
     X"a9", X"10", X"85", X"99", X"a2", X"00", X"a0", X"00",
     X"8a", X"0a", X"aa", X"98", X"2a", X"a8", X"b0", X"a4",
     X"06", X"ad", X"26", X"ae", X"90", X"0b", X"18", X"8a",
     X"65", X"64", X"aa", X"98", X"65", X"65", X"a8", X"b0",
     X"93", X"c6", X"99", X"d0", X"e3", X"60", X"a5", X"11",
     X"f0", X"03", X"20", X"00", X"e6", X"20", X"84", X"e4",
     X"38", X"a5", X"6f", X"e5", X"6d", X"a8", X"a5", X"70",
     X"e5", X"6e", X"a2", X"00", X"86", X"11", X"85", X"9e",
     X"84", X"9f", X"a2", X"90", X"4c", X"9b", X"eb", X"a4",
     X"24", X"a9", X"00", X"38", X"f0", X"ec", X"a6", X"76",
     X"e8", X"d0", X"a1", X"a2", X"95", X"2c", X"a2", X"e0",
     X"4c", X"12", X"d4", X"20", X"41", X"e3", X"20", X"06",
     X"e3", X"20", X"bb", X"de", X"a9", X"80", X"85", X"14",
     X"20", X"e3", X"df", X"20", X"6a", X"dd", X"20", X"b8",
     X"de", X"a9", X"d0", X"20", X"c0", X"de", X"48", X"a5",
     X"84", X"48", X"a5", X"83", X"48", X"a5", X"b9", X"48",
     X"a5", X"b8", X"48", X"20", X"95", X"d9", X"4c", X"af",
     X"e3", X"a9", X"c2", X"20", X"c0", X"de", X"09", X"80",
     X"85", X"14", X"20", X"ea", X"df", X"85", X"8a", X"84",
     X"8b", X"4c", X"6a", X"dd", X"20", X"41", X"e3", X"a5",
     X"8b", X"48", X"a5", X"8a", X"48", X"20", X"b2", X"de",
     X"20", X"6a", X"dd", X"68", X"85", X"8a", X"68", X"85",
     X"8b", X"a0", X"02", X"b1", X"8a", X"85", X"83", X"aa",
     X"c8", X"b1", X"8a", X"f0", X"99", X"85", X"84", X"c8",
     X"b1", X"83", X"48", X"88", X"10", X"fa", X"a4", X"84",
     X"20", X"2b", X"eb", X"a5", X"b9", X"48", X"a5", X"b8",
     X"48", X"b1", X"8a", X"85", X"b8", X"c8", X"b1", X"8a",
     X"85", X"b9", X"a5", X"84", X"48", X"a5", X"83", X"48",
     X"20", X"67", X"dd", X"68", X"85", X"8a", X"68", X"85",
     X"8b", X"20", X"b7", X"00", X"f0", X"03", X"4c", X"c9",
     X"de", X"68", X"85", X"b8", X"68", X"85", X"b9", X"a0",
     X"00", X"68", X"91", X"8a", X"68", X"c8", X"91", X"8a",
     X"68", X"c8", X"91", X"8a", X"68", X"c8", X"91", X"8a",
     X"68", X"c8", X"91", X"8a", X"60", X"20", X"6a", X"dd",
     X"a0", X"00", X"20", X"36", X"ed", X"68", X"68", X"a9",
     X"ff", X"a0", X"00", X"f0", X"12", X"a6", X"a0", X"a4",
     X"a1", X"86", X"8c", X"84", X"8d", X"20", X"52", X"e4",
     X"86", X"9e", X"84", X"9f", X"85", X"9d", X"60", X"a2",
     X"22", X"86", X"0d", X"86", X"0e", X"85", X"ab", X"84",
     X"ac", X"85", X"9e", X"84", X"9f", X"a0", X"ff", X"c8",
     X"b1", X"ab", X"f0", X"0c", X"c5", X"0d", X"f0", X"04",
     X"c5", X"0e", X"d0", X"f3", X"c9", X"22", X"f0", X"01",
     X"18", X"84", X"9d", X"98", X"65", X"ab", X"85", X"ad",
     X"a6", X"ac", X"90", X"01", X"e8", X"86", X"ae", X"a5",
     X"ac", X"f0", X"04", X"c9", X"02", X"d0", X"0b", X"98",
     X"20", X"d5", X"e3", X"a6", X"ab", X"a4", X"ac", X"20",
     X"e2", X"e5", X"a6", X"52", X"e0", X"5e", X"d0", X"05",
     X"a2", X"bf", X"4c", X"12", X"d4", X"a5", X"9d", X"95",
     X"00", X"a5", X"9e", X"95", X"01", X"a5", X"9f", X"95",
     X"02", X"a0", X"00", X"86", X"a0", X"84", X"a1", X"88",
     X"84", X"11", X"86", X"53", X"e8", X"e8", X"e8", X"86",
     X"52", X"60", X"46", X"13", X"48", X"49", X"ff", X"38",
     X"65", X"6f", X"a4", X"70", X"b0", X"01", X"88", X"c4",
     X"6e", X"90", X"11", X"d0", X"04", X"c5", X"6d", X"90",
     X"0b", X"85", X"6f", X"84", X"70", X"85", X"71", X"84",
     X"72", X"aa", X"68", X"60", X"a2", X"4d", X"a5", X"13",
     X"30", X"b8", X"20", X"84", X"e4", X"a9", X"80", X"85",
     X"13", X"68", X"d0", X"d0", X"a6", X"73", X"a5", X"74",
     X"86", X"6f", X"85", X"70", X"a0", X"00", X"84", X"8b",
     X"a5", X"6d", X"a6", X"6e", X"85", X"9b", X"86", X"9c",
     X"a9", X"55", X"a2", X"00", X"85", X"5e", X"86", X"5f",
     X"c5", X"52", X"f0", X"05", X"20", X"23", X"e5", X"f0",
     X"f7", X"a9", X"07", X"85", X"8f", X"a5", X"69", X"a6",
     X"6a", X"85", X"5e", X"86", X"5f", X"e4", X"6c", X"d0",
     X"04", X"c5", X"6b", X"f0", X"05", X"20", X"19", X"e5",
     X"f0", X"f3", X"85", X"94", X"86", X"95", X"a9", X"03",
     X"85", X"8f", X"a5", X"94", X"a6", X"95", X"e4", X"6e",
     X"d0", X"07", X"c5", X"6d", X"d0", X"03", X"4c", X"62",
     X"e5", X"85", X"5e", X"86", X"5f", X"a0", X"00", X"b1",
     X"5e", X"aa", X"c8", X"b1", X"5e", X"08", X"c8", X"b1",
     X"5e", X"65", X"94", X"85", X"94", X"c8", X"b1", X"5e",
     X"65", X"95", X"85", X"95", X"28", X"10", X"d3", X"8a",
     X"30", X"d0", X"c8", X"b1", X"5e", X"a0", X"00", X"0a",
     X"69", X"05", X"65", X"5e", X"85", X"5e", X"90", X"02",
     X"e6", X"5f", X"a6", X"5f", X"e4", X"95", X"d0", X"04",
     X"c5", X"94", X"f0", X"ba", X"20", X"23", X"e5", X"f0",
     X"f3", X"b1", X"5e", X"30", X"35", X"c8", X"b1", X"5e",
     X"10", X"30", X"c8", X"b1", X"5e", X"f0", X"2b", X"c8",
     X"b1", X"5e", X"aa", X"c8", X"b1", X"5e", X"c5", X"70",
     X"90", X"06", X"d0", X"1e", X"e4", X"6f", X"b0", X"1a",
     X"c5", X"9c", X"90", X"16", X"d0", X"04", X"e4", X"9b",
     X"90", X"10", X"86", X"9b", X"85", X"9c", X"a5", X"5e",
     X"a6", X"5f", X"85", X"8a", X"86", X"8b", X"a5", X"8f",
     X"85", X"91", X"a5", X"8f", X"18", X"65", X"5e", X"85",
     X"5e", X"90", X"02", X"e6", X"5f", X"a6", X"5f", X"a0",
     X"00", X"60", X"a6", X"8b", X"f0", X"f7", X"a5", X"91",
     X"29", X"04", X"4a", X"a8", X"85", X"91", X"b1", X"8a",
     X"65", X"9b", X"85", X"96", X"a5", X"9c", X"69", X"00",
     X"85", X"97", X"a5", X"6f", X"a6", X"70", X"85", X"94",
     X"86", X"95", X"20", X"9a", X"d3", X"a4", X"91", X"c8",
     X"a5", X"94", X"91", X"8a", X"aa", X"e6", X"95", X"a5",
     X"95", X"c8", X"91", X"8a", X"4c", X"88", X"e4", X"a5",
     X"a1", X"48", X"a5", X"a0", X"48", X"20", X"60", X"de",
     X"20", X"6c", X"dd", X"68", X"85", X"ab", X"68", X"85",
     X"ac", X"a0", X"00", X"b1", X"ab", X"18", X"71", X"a0",
     X"90", X"05", X"a2", X"b0", X"4c", X"12", X"d4", X"20",
     X"d5", X"e3", X"20", X"d4", X"e5", X"a5", X"8c", X"a4",
     X"8d", X"20", X"04", X"e6", X"20", X"e6", X"e5", X"a5",
     X"ab", X"a4", X"ac", X"20", X"04", X"e6", X"20", X"2a",
     X"e4", X"4c", X"95", X"dd", X"a0", X"00", X"b1", X"ab",
     X"48", X"c8", X"b1", X"ab", X"aa", X"c8", X"b1", X"ab",
     X"a8", X"68", X"86", X"5e", X"84", X"5f", X"a8", X"f0",
     X"0a", X"48", X"88", X"b1", X"5e", X"91", X"71", X"98",
     X"d0", X"f8", X"68", X"18", X"65", X"71", X"85", X"71",
     X"90", X"02", X"e6", X"72", X"60", X"20", X"6c", X"dd",
     X"a5", X"a0", X"a4", X"a1", X"85", X"5e", X"84", X"5f",
     X"20", X"35", X"e6", X"08", X"a0", X"00", X"b1", X"5e",
     X"48", X"c8", X"b1", X"5e", X"aa", X"c8", X"b1", X"5e",
     X"a8", X"68", X"28", X"d0", X"13", X"c4", X"70", X"d0",
     X"0f", X"e4", X"6f", X"d0", X"0b", X"48", X"18", X"65",
     X"6f", X"85", X"6f", X"90", X"02", X"e6", X"70", X"68",
     X"86", X"5e", X"84", X"5f", X"60", X"c4", X"54", X"d0",
     X"0c", X"c5", X"53", X"d0", X"08", X"85", X"52", X"e9",
     X"03", X"85", X"53", X"a0", X"00", X"60", X"20", X"fb",
     X"e6", X"8a", X"48", X"a9", X"01", X"20", X"dd", X"e3",
     X"68", X"a0", X"00", X"91", X"9e", X"68", X"68", X"4c",
     X"2a", X"e4", X"20", X"b9", X"e6", X"d1", X"8c", X"98",
     X"90", X"04", X"b1", X"8c", X"aa", X"98", X"48", X"8a",
     X"48", X"20", X"dd", X"e3", X"a5", X"8c", X"a4", X"8d",
     X"20", X"04", X"e6", X"68", X"a8", X"68", X"18", X"65",
     X"5e", X"85", X"5e", X"90", X"02", X"e6", X"5f", X"98",
     X"20", X"e6", X"e5", X"4c", X"2a", X"e4", X"20", X"b9",
     X"e6", X"18", X"f1", X"8c", X"49", X"ff", X"4c", X"60",
     X"e6", X"a9", X"ff", X"85", X"a1", X"20", X"b7", X"00",
     X"c9", X"29", X"f0", X"06", X"20", X"be", X"de", X"20",
     X"f8", X"e6", X"20", X"b9", X"e6", X"ca", X"8a", X"48",
     X"18", X"a2", X"00", X"f1", X"8c", X"b0", X"b8", X"49",
     X"ff", X"c5", X"a1", X"90", X"b3", X"a5", X"a1", X"b0",
     X"af", X"20", X"b8", X"de", X"68", X"a8", X"68", X"85",
     X"91", X"68", X"68", X"68", X"aa", X"68", X"85", X"8c",
     X"68", X"85", X"8d", X"a5", X"91", X"48", X"98", X"48",
     X"a0", X"00", X"8a", X"f0", X"1d", X"60", X"20", X"dc",
     X"e6", X"4c", X"01", X"e3", X"20", X"fd", X"e5", X"a2",
     X"00", X"86", X"11", X"a8", X"60", X"20", X"dc", X"e6",
     X"f0", X"08", X"a0", X"00", X"b1", X"5e", X"a8", X"4c",
     X"01", X"e3", X"4c", X"99", X"e1", X"20", X"b1", X"00",
     X"20", X"67", X"dd", X"20", X"08", X"e1", X"a6", X"a0",
     X"d0", X"f0", X"a6", X"a1", X"4c", X"b7", X"00", X"20",
     X"dc", X"e6", X"d0", X"03", X"4c", X"4e", X"e8", X"a6",
     X"b8", X"a4", X"b9", X"86", X"ad", X"84", X"ae", X"a6",
     X"5e", X"86", X"b8", X"18", X"65", X"5e", X"85", X"60",
     X"a6", X"5f", X"86", X"b9", X"90", X"01", X"e8", X"86",
     X"61", X"a0", X"00", X"b1", X"60", X"48", X"a9", X"00",
     X"91", X"60", X"20", X"b7", X"00", X"20", X"4a", X"ec",
     X"68", X"a0", X"00", X"91", X"60", X"a6", X"ad", X"a4",
     X"ae", X"86", X"b8", X"84", X"b9", X"60", X"20", X"67",
     X"dd", X"20", X"52", X"e7", X"20", X"be", X"de", X"4c",
     X"f8", X"e6", X"a5", X"9d", X"c9", X"91", X"b0", X"9a",
     X"20", X"f2", X"eb", X"a5", X"a0", X"a4", X"a1", X"84",
     X"50", X"85", X"51", X"60", X"a5", X"50", X"48", X"a5",
     X"51", X"48", X"20", X"52", X"e7", X"a0", X"00", X"b1",
     X"50", X"a8", X"68", X"85", X"51", X"68", X"85", X"50",
     X"4c", X"01", X"e3", X"20", X"46", X"e7", X"8a", X"a0",
     X"00", X"91", X"50", X"60", X"20", X"46", X"e7", X"86",
     X"85", X"a2", X"00", X"20", X"b7", X"00", X"f0", X"03",
     X"20", X"4c", X"e7", X"86", X"86", X"a0", X"00", X"b1",
     X"50", X"45", X"86", X"25", X"85", X"f0", X"f8", X"60",
     X"a9", X"64", X"a0", X"ee", X"4c", X"be", X"e7", X"20",
     X"e3", X"e9", X"a5", X"a2", X"49", X"ff", X"85", X"a2",
     X"45", X"aa", X"85", X"ab", X"a5", X"9d", X"4c", X"c1",
     X"e7", X"20", X"f0", X"e8", X"90", X"3c", X"20", X"e3",
     X"e9", X"d0", X"03", X"4c", X"53", X"eb", X"a6", X"ac",
     X"86", X"92", X"a2", X"a5", X"a5", X"a5", X"a8", X"f0",
     X"ce", X"38", X"e5", X"9d", X"f0", X"24", X"90", X"12",
     X"84", X"9d", X"a4", X"aa", X"84", X"a2", X"49", X"ff",
     X"69", X"00", X"a0", X"00", X"84", X"92", X"a2", X"9d",
     X"d0", X"04", X"a0", X"00", X"84", X"ac", X"c9", X"f9",
     X"30", X"c7", X"a8", X"a5", X"ac", X"56", X"01", X"20",
     X"07", X"e9", X"24", X"ab", X"10", X"57", X"a0", X"9d",
     X"e0", X"a5", X"f0", X"02", X"a0", X"a5", X"38", X"49",
     X"ff", X"65", X"92", X"85", X"ac", X"b9", X"04", X"00",
     X"f5", X"04", X"85", X"a1", X"b9", X"03", X"00", X"f5",
     X"03", X"85", X"a0", X"b9", X"02", X"00", X"f5", X"02",
     X"85", X"9f", X"b9", X"01", X"00", X"f5", X"01", X"85",
     X"9e", X"b0", X"03", X"20", X"9e", X"e8", X"a0", X"00",
     X"98", X"18", X"a6", X"9e", X"d0", X"4a", X"a6", X"9f",
     X"86", X"9e", X"a6", X"a0", X"86", X"9f", X"a6", X"a1",
     X"86", X"a0", X"a6", X"ac", X"86", X"a1", X"84", X"ac",
     X"69", X"08", X"c9", X"20", X"d0", X"e4", X"a9", X"00",
     X"85", X"9d", X"85", X"a2", X"60", X"65", X"92", X"85",
     X"ac", X"a5", X"a1", X"65", X"a9", X"85", X"a1", X"a5",
     X"a0", X"65", X"a8", X"85", X"a0", X"a5", X"9f", X"65",
     X"a7", X"85", X"9f", X"a5", X"9e", X"65", X"a6", X"85",
     X"9e", X"4c", X"8d", X"e8", X"69", X"01", X"06", X"ac",
     X"26", X"a1", X"26", X"a0", X"26", X"9f", X"26", X"9e",
     X"10", X"f2", X"38", X"e5", X"9d", X"b0", X"c7", X"49",
     X"ff", X"69", X"01", X"85", X"9d", X"90", X"0e", X"e6",
     X"9d", X"f0", X"42", X"66", X"9e", X"66", X"9f", X"66",
     X"a0", X"66", X"a1", X"66", X"ac", X"60", X"a5", X"a2",
     X"49", X"ff", X"85", X"a2", X"a5", X"9e", X"49", X"ff",
     X"85", X"9e", X"a5", X"9f", X"49", X"ff", X"85", X"9f",
     X"a5", X"a0", X"49", X"ff", X"85", X"a0", X"a5", X"a1",
     X"49", X"ff", X"85", X"a1", X"a5", X"ac", X"49", X"ff",
     X"85", X"ac", X"e6", X"ac", X"d0", X"0e", X"e6", X"a1",
     X"d0", X"0a", X"e6", X"a0", X"d0", X"06", X"e6", X"9f",
     X"d0", X"02", X"e6", X"9e", X"60", X"a2", X"45", X"4c",
     X"12", X"d4", X"a2", X"61", X"b4", X"04", X"84", X"ac",
     X"b4", X"03", X"94", X"04", X"b4", X"02", X"94", X"03",
     X"b4", X"01", X"94", X"02", X"a4", X"a4", X"94", X"01",
     X"69", X"08", X"30", X"e8", X"f0", X"e6", X"e9", X"08",
     X"a8", X"a5", X"ac", X"b0", X"14", X"16", X"01", X"90",
     X"02", X"f6", X"01", X"76", X"01", X"76", X"01", X"76",
     X"02", X"76", X"03", X"76", X"04", X"6a", X"c8", X"d0",
     X"ec", X"18", X"60", X"81", X"00", X"00", X"00", X"00",
     X"03", X"7f", X"5e", X"56", X"cb", X"79", X"80", X"13",
     X"9b", X"0b", X"64", X"80", X"76", X"38", X"93", X"16",
     X"82", X"38", X"aa", X"3b", X"20", X"80", X"35", X"04",
     X"f3", X"34", X"81", X"35", X"04", X"f3", X"34", X"80",
     X"80", X"00", X"00", X"00", X"80", X"31", X"72", X"17",
     X"f8", X"20", X"82", X"eb", X"f0", X"02", X"10", X"03",
     X"4c", X"99", X"e1", X"a5", X"9d", X"e9", X"7f", X"48",
     X"a9", X"80", X"85", X"9d", X"a9", X"2d", X"a0", X"e9",
     X"20", X"be", X"e7", X"a9", X"32", X"a0", X"e9", X"20",
     X"66", X"ea", X"a9", X"13", X"a0", X"e9", X"20", X"a7",
     X"e7", X"a9", X"18", X"a0", X"e9", X"20", X"5c", X"ef",
     X"a9", X"37", X"a0", X"e9", X"20", X"be", X"e7", X"68",
     X"20", X"d5", X"ec", X"a9", X"3c", X"a0", X"e9", X"20",
     X"e3", X"e9", X"d0", X"03", X"4c", X"e2", X"e9", X"20",
     X"0e", X"ea", X"a9", X"00", X"85", X"62", X"85", X"63",
     X"85", X"64", X"85", X"65", X"a5", X"ac", X"20", X"b0",
     X"e9", X"a5", X"a1", X"20", X"b0", X"e9", X"a5", X"a0",
     X"20", X"b0", X"e9", X"a5", X"9f", X"20", X"b0", X"e9",
     X"a5", X"9e", X"20", X"b5", X"e9", X"4c", X"e6", X"ea",
     X"d0", X"03", X"4c", X"da", X"e8", X"4a", X"09", X"80",
     X"a8", X"90", X"19", X"18", X"a5", X"65", X"65", X"a9",
     X"85", X"65", X"a5", X"64", X"65", X"a8", X"85", X"64",
     X"a5", X"63", X"65", X"a7", X"85", X"63", X"a5", X"62",
     X"65", X"a6", X"85", X"62", X"66", X"62", X"66", X"63",
     X"66", X"64", X"66", X"65", X"66", X"ac", X"98", X"4a",
     X"d0", X"d6", X"60", X"85", X"5e", X"84", X"5f", X"a0",
     X"04", X"b1", X"5e", X"85", X"a9", X"88", X"b1", X"5e",
     X"85", X"a8", X"88", X"b1", X"5e", X"85", X"a7", X"88",
     X"b1", X"5e", X"85", X"aa", X"45", X"a2", X"85", X"ab",
     X"a5", X"aa", X"09", X"80", X"85", X"a6", X"88", X"b1",
     X"5e", X"85", X"a5", X"a5", X"9d", X"60", X"a5", X"a5",
     X"f0", X"1f", X"18", X"65", X"9d", X"90", X"04", X"30",
     X"1d", X"18", X"2c", X"10", X"14", X"69", X"80", X"85",
     X"9d", X"d0", X"03", X"4c", X"52", X"e8", X"a5", X"ab",
     X"85", X"a2", X"60", X"a5", X"a2", X"49", X"ff", X"30",
     X"05", X"68", X"68", X"4c", X"4e", X"e8", X"4c", X"d5",
     X"e8", X"20", X"63", X"eb", X"aa", X"f0", X"10", X"18",
     X"69", X"02", X"b0", X"f2", X"a2", X"00", X"86", X"ab",
     X"20", X"ce", X"e7", X"e6", X"9d", X"f0", X"e7", X"60",
     X"84", X"20", X"00", X"00", X"00", X"20", X"63", X"eb",
     X"a9", X"50", X"a0", X"ea", X"a2", X"00", X"86", X"ab",
     X"20", X"f9", X"ea", X"4c", X"69", X"ea", X"20", X"e3",
     X"e9", X"f0", X"76", X"20", X"72", X"eb", X"a9", X"00",
     X"38", X"e5", X"9d", X"85", X"9d", X"20", X"0e", X"ea",
     X"e6", X"9d", X"f0", X"ba", X"a2", X"fc", X"a9", X"01",
     X"a4", X"a6", X"c4", X"9e", X"d0", X"10", X"a4", X"a7",
     X"c4", X"9f", X"d0", X"0a", X"a4", X"a8", X"c4", X"a0",
     X"d0", X"04", X"a4", X"a9", X"c4", X"a1", X"08", X"2a",
     X"90", X"09", X"e8", X"95", X"65", X"f0", X"32", X"10",
     X"34", X"a9", X"01", X"28", X"b0", X"0e", X"06", X"a9",
     X"26", X"a8", X"26", X"a7", X"26", X"a6", X"b0", X"e6",
     X"30", X"ce", X"10", X"e2", X"a8", X"a5", X"a9", X"e5",
     X"a1", X"85", X"a9", X"a5", X"a8", X"e5", X"a0", X"85",
     X"a8", X"a5", X"a7", X"e5", X"9f", X"85", X"a7", X"a5",
     X"a6", X"e5", X"9e", X"85", X"a6", X"98", X"4c", X"a6",
     X"ea", X"a9", X"40", X"d0", X"ce", X"0a", X"0a", X"0a",
     X"0a", X"0a", X"0a", X"85", X"ac", X"28", X"4c", X"e6",
     X"ea", X"a2", X"85", X"4c", X"12", X"d4", X"a5", X"62",
     X"85", X"9e", X"a5", X"63", X"85", X"9f", X"a5", X"64",
     X"85", X"a0", X"a5", X"65", X"85", X"a1", X"4c", X"2e",
     X"e8", X"85", X"5e", X"84", X"5f", X"a0", X"04", X"b1",
     X"5e", X"85", X"a1", X"88", X"b1", X"5e", X"85", X"a0",
     X"88", X"b1", X"5e", X"85", X"9f", X"88", X"b1", X"5e",
     X"85", X"a2", X"09", X"80", X"85", X"9e", X"88", X"b1",
     X"5e", X"85", X"9d", X"84", X"ac", X"60", X"a2", X"98",
     X"2c", X"a2", X"93", X"a0", X"00", X"f0", X"04", X"a6",
     X"85", X"a4", X"86", X"20", X"72", X"eb", X"86", X"5e",
     X"84", X"5f", X"a0", X"04", X"a5", X"a1", X"91", X"5e",
     X"88", X"a5", X"a0", X"91", X"5e", X"88", X"a5", X"9f",
     X"91", X"5e", X"88", X"a5", X"a2", X"09", X"7f", X"25",
     X"9e", X"91", X"5e", X"88", X"a5", X"9d", X"91", X"5e",
     X"84", X"ac", X"60", X"a5", X"aa", X"85", X"a2", X"a2",
     X"05", X"b5", X"a4", X"95", X"9c", X"ca", X"d0", X"f9",
     X"86", X"ac", X"60", X"20", X"72", X"eb", X"a2", X"06",
     X"b5", X"9c", X"95", X"a4", X"ca", X"d0", X"f9", X"86",
     X"ac", X"60", X"a5", X"9d", X"f0", X"fb", X"06", X"ac",
     X"90", X"f7", X"20", X"c6", X"e8", X"d0", X"f2", X"4c",
     X"8f", X"e8", X"a5", X"9d", X"f0", X"09", X"a5", X"a2",
     X"2a", X"a9", X"ff", X"b0", X"02", X"a9", X"01", X"60",
     X"20", X"82", X"eb", X"85", X"9e", X"a9", X"00", X"85",
     X"9f", X"a2", X"88", X"a5", X"9e", X"49", X"ff", X"2a",
     X"a9", X"00", X"85", X"a1", X"85", X"a0", X"86", X"9d",
     X"85", X"ac", X"85", X"a2", X"4c", X"29", X"e8", X"46",
     X"a2", X"60", X"85", X"60", X"84", X"61", X"a0", X"00",
     X"b1", X"60", X"c8", X"aa", X"f0", X"c4", X"b1", X"60",
     X"45", X"a2", X"30", X"c2", X"e4", X"9d", X"d0", X"21",
     X"b1", X"60", X"09", X"80", X"c5", X"9e", X"d0", X"19",
     X"c8", X"b1", X"60", X"c5", X"9f", X"d0", X"12", X"c8",
     X"b1", X"60", X"c5", X"a0", X"d0", X"0b", X"c8", X"a9",
     X"7f", X"c5", X"ac", X"b1", X"60", X"e5", X"a1", X"f0",
     X"28", X"a5", X"a2", X"90", X"02", X"49", X"ff", X"4c",
     X"88", X"eb", X"a5", X"9d", X"f0", X"4a", X"38", X"e9",
     X"a0", X"24", X"a2", X"10", X"09", X"aa", X"a9", X"ff",
     X"85", X"a4", X"20", X"a4", X"e8", X"8a", X"a2", X"9d",
     X"c9", X"f9", X"10", X"06", X"20", X"f0", X"e8", X"84",
     X"a4", X"60", X"a8", X"a5", X"a2", X"29", X"80", X"46",
     X"9e", X"05", X"9e", X"85", X"9e", X"20", X"07", X"e9",
     X"84", X"a4", X"60", X"a5", X"9d", X"c9", X"a0", X"b0",
     X"20", X"20", X"f2", X"eb", X"84", X"ac", X"a5", X"a2",
     X"84", X"a2", X"49", X"80", X"2a", X"a9", X"a0", X"85",
     X"9d", X"a5", X"a1", X"85", X"0d", X"4c", X"29", X"e8",
     X"85", X"9e", X"85", X"9f", X"85", X"a0", X"85", X"a1",
     X"a8", X"60", X"a0", X"00", X"a2", X"0a", X"94", X"99",
     X"ca", X"10", X"fb", X"90", X"0f", X"c9", X"2d", X"d0",
     X"04", X"86", X"a3", X"f0", X"04", X"c9", X"2b", X"d0",
     X"05", X"20", X"b1", X"00", X"90", X"5b", X"c9", X"2e",
     X"f0", X"2e", X"c9", X"45", X"d0", X"30", X"20", X"b1",
     X"00", X"90", X"17", X"c9", X"c9", X"f0", X"0e", X"c9",
     X"2d", X"f0", X"0a", X"c9", X"c8", X"f0", X"08", X"c9",
     X"2b", X"f0", X"04", X"d0", X"07", X"66", X"9c", X"20",
     X"b1", X"00", X"90", X"5c", X"24", X"9c", X"10", X"0e",
     X"a9", X"00", X"38", X"e5", X"9a", X"4c", X"a0", X"ec",
     X"66", X"9b", X"24", X"9b", X"50", X"c3", X"a5", X"9a",
     X"38", X"e5", X"99", X"85", X"9a", X"f0", X"12", X"10",
     X"09", X"20", X"55", X"ea", X"e6", X"9a", X"d0", X"f9",
     X"f0", X"07", X"20", X"39", X"ea", X"c6", X"9a", X"d0",
     X"f9", X"a5", X"a3", X"30", X"01", X"60", X"4c", X"d0",
     X"ee", X"48", X"24", X"9b", X"10", X"02", X"e6", X"99",
     X"20", X"39", X"ea", X"68", X"38", X"e9", X"30", X"20",
     X"d5", X"ec", X"4c", X"61", X"ec", X"48", X"20", X"63",
     X"eb", X"68", X"20", X"93", X"eb", X"a5", X"aa", X"45",
     X"a2", X"85", X"ab", X"a6", X"9d", X"4c", X"c1", X"e7",
     X"a5", X"9a", X"c9", X"0a", X"90", X"09", X"a9", X"64",
     X"24", X"9c", X"30", X"11", X"4c", X"d5", X"e8", X"0a",
     X"0a", X"18", X"65", X"9a", X"0a", X"18", X"a0", X"00",
     X"71", X"b8", X"38", X"e9", X"30", X"85", X"9a", X"4c",
     X"87", X"ec", X"9b", X"3e", X"bc", X"1f", X"fd", X"9e",
     X"6e", X"6b", X"27", X"fd", X"9e", X"6e", X"6b", X"28",
     X"00", X"a9", X"58", X"a0", X"d3", X"20", X"31", X"ed",
     X"a5", X"76", X"a6", X"75", X"85", X"9e", X"86", X"9f",
     X"a2", X"90", X"38", X"20", X"a0", X"eb", X"20", X"34",
     X"ed", X"4c", X"3a", X"db", X"a0", X"01", X"a9", X"2d",
     X"88", X"24", X"a2", X"10", X"04", X"c8", X"99", X"ff",
     X"00", X"85", X"a2", X"84", X"ad", X"c8", X"a9", X"30",
     X"a6", X"9d", X"d0", X"03", X"4c", X"57", X"ee", X"a9",
     X"00", X"e0", X"80", X"f0", X"02", X"b0", X"09", X"a9",
     X"14", X"a0", X"ed", X"20", X"7f", X"e9", X"a9", X"f7",
     X"85", X"99", X"a9", X"0f", X"a0", X"ed", X"20", X"b2",
     X"eb", X"f0", X"1e", X"10", X"12", X"a9", X"0a", X"a0",
     X"ed", X"20", X"b2", X"eb", X"f0", X"02", X"10", X"0e",
     X"20", X"39", X"ea", X"c6", X"99", X"d0", X"ee", X"20",
     X"55", X"ea", X"e6", X"99", X"d0", X"dc", X"20", X"a0",
     X"e7", X"20", X"f2", X"eb", X"a2", X"01", X"a5", X"99",
     X"18", X"69", X"0a", X"30", X"09", X"c9", X"0b", X"b0",
     X"06", X"69", X"ff", X"aa", X"a9", X"02", X"38", X"e9",
     X"02", X"85", X"9a", X"86", X"99", X"8a", X"f0", X"02",
     X"10", X"13", X"a4", X"ad", X"a9", X"2e", X"c8", X"99",
     X"ff", X"00", X"8a", X"f0", X"06", X"a9", X"30", X"c8",
     X"99", X"ff", X"00", X"84", X"ad", X"a0", X"00", X"a2",
     X"80", X"a5", X"a1", X"18", X"79", X"6c", X"ee", X"85",
     X"a1", X"a5", X"a0", X"79", X"6b", X"ee", X"85", X"a0",
     X"a5", X"9f", X"79", X"6a", X"ee", X"85", X"9f", X"a5",
     X"9e", X"79", X"69", X"ee", X"85", X"9e", X"e8", X"b0",
     X"04", X"10", X"de", X"30", X"02", X"30", X"da", X"8a",
     X"90", X"04", X"49", X"ff", X"69", X"0a", X"69", X"2f",
     X"c8", X"c8", X"c8", X"c8", X"84", X"83", X"a4", X"ad",
     X"c8", X"aa", X"29", X"7f", X"99", X"ff", X"00", X"c6",
     X"99", X"d0", X"06", X"a9", X"2e", X"c8", X"99", X"ff",
     X"00", X"84", X"ad", X"a4", X"83", X"8a", X"49", X"ff",
     X"29", X"80", X"aa", X"c0", X"24", X"d0", X"aa", X"a4",
     X"ad", X"b9", X"ff", X"00", X"88", X"c9", X"30", X"f0",
     X"f8", X"c9", X"2e", X"f0", X"01", X"c8", X"a9", X"2b",
     X"a6", X"9a", X"f0", X"2e", X"10", X"08", X"a9", X"00",
     X"38", X"e5", X"9a", X"aa", X"a9", X"2d", X"99", X"01",
     X"01", X"a9", X"45", X"99", X"00", X"01", X"8a", X"a2",
     X"2f", X"38", X"e8", X"e9", X"0a", X"b0", X"fb", X"69",
     X"3a", X"99", X"03", X"01", X"8a", X"99", X"02", X"01",
     X"a9", X"00", X"99", X"04", X"01", X"f0", X"08", X"99",
     X"ff", X"00", X"a9", X"00", X"99", X"00", X"01", X"a9",
     X"00", X"a0", X"01", X"60", X"80", X"00", X"00", X"00",
     X"00", X"fa", X"0a", X"1f", X"00", X"00", X"98", X"96",
     X"80", X"ff", X"f0", X"bd", X"c0", X"00", X"01", X"86",
     X"a0", X"ff", X"ff", X"d8", X"f0", X"00", X"00", X"03",
     X"e8", X"ff", X"ff", X"ff", X"9c", X"00", X"00", X"00",
     X"0a", X"ff", X"ff", X"ff", X"ff", X"20", X"63", X"eb",
     X"a9", X"64", X"a0", X"ee", X"20", X"f9", X"ea", X"f0",
     X"70", X"a5", X"a5", X"d0", X"03", X"4c", X"50", X"e8",
     X"a2", X"8a", X"a0", X"00", X"20", X"2b", X"eb", X"a5",
     X"aa", X"10", X"0f", X"20", X"23", X"ec", X"a9", X"8a",
     X"a0", X"00", X"20", X"b2", X"eb", X"d0", X"03", X"98",
     X"a4", X"0d", X"20", X"55", X"eb", X"98", X"48", X"20",
     X"41", X"e9", X"a9", X"8a", X"a0", X"00", X"20", X"7f",
     X"e9", X"20", X"09", X"ef", X"68", X"4a", X"90", X"0a",
     X"a5", X"9d", X"f0", X"06", X"a5", X"a2", X"49", X"ff",
     X"85", X"a2", X"60", X"81", X"38", X"aa", X"3b", X"29",
     X"07", X"71", X"34", X"58", X"3e", X"56", X"74", X"16",
     X"7e", X"b3", X"1b", X"77", X"2f", X"ee", X"e3", X"85",
     X"7a", X"1d", X"84", X"1c", X"2a", X"7c", X"63", X"59",
     X"58", X"0a", X"7e", X"75", X"fd", X"e7", X"c6", X"80",
     X"31", X"72", X"18", X"10", X"81", X"00", X"00", X"00",
     X"00", X"a9", X"db", X"a0", X"ee", X"20", X"7f", X"e9",
     X"a5", X"ac", X"69", X"50", X"90", X"03", X"20", X"7a",
     X"eb", X"85", X"92", X"20", X"66", X"eb", X"a5", X"9d",
     X"c9", X"88", X"90", X"03", X"20", X"2b", X"ea", X"20",
     X"23", X"ec", X"a5", X"0d", X"18", X"69", X"81", X"f0",
     X"f3", X"38", X"e9", X"01", X"48", X"a2", X"05", X"b5",
     X"a5", X"b4", X"9d", X"95", X"9d", X"94", X"a5", X"ca",
     X"10", X"f5", X"a5", X"92", X"85", X"ac", X"20", X"aa",
     X"e7", X"20", X"d0", X"ee", X"a9", X"e0", X"a0", X"ee",
     X"20", X"72", X"ef", X"a9", X"00", X"85", X"ab", X"68",
     X"20", X"10", X"ea", X"60", X"85", X"ad", X"84", X"ae",
     X"20", X"21", X"eb", X"a9", X"93", X"20", X"7f", X"e9",
     X"20", X"76", X"ef", X"a9", X"93", X"a0", X"00", X"4c",
     X"7f", X"e9", X"85", X"ad", X"84", X"ae", X"20", X"1e",
     X"eb", X"b1", X"ad", X"85", X"a3", X"a4", X"ad", X"c8",
     X"98", X"d0", X"02", X"e6", X"ae", X"85", X"ad", X"a4",
     X"ae", X"20", X"7f", X"e9", X"a5", X"ad", X"a4", X"ae",
     X"18", X"69", X"05", X"90", X"01", X"c8", X"85", X"ad",
     X"84", X"ae", X"20", X"be", X"e7", X"a9", X"98", X"a0",
     X"00", X"c6", X"a3", X"d0", X"e4", X"60", X"98", X"35",
     X"44", X"7a", X"68", X"28", X"b1", X"46", X"20", X"82",
     X"eb", X"aa", X"30", X"18", X"a9", X"c9", X"a0", X"00",
     X"20", X"f9", X"ea", X"8a", X"f0", X"e7", X"a9", X"a6",
     X"a0", X"ef", X"20", X"7f", X"e9", X"a9", X"aa", X"a0",
     X"ef", X"20", X"be", X"e7", X"a6", X"a1", X"a5", X"9e",
     X"85", X"a1", X"86", X"9e", X"a9", X"00", X"85", X"a2",
     X"a5", X"9d", X"85", X"ac", X"a9", X"80", X"85", X"9d",
     X"20", X"2e", X"e8", X"a2", X"c9", X"a0", X"00", X"4c",
     X"2b", X"eb", X"a9", X"66", X"a0", X"f0", X"20", X"be",
     X"e7", X"20", X"63", X"eb", X"a9", X"6b", X"a0", X"f0",
     X"a6", X"aa", X"20", X"5e", X"ea", X"20", X"63", X"eb",
     X"20", X"23", X"ec", X"a9", X"00", X"85", X"ab", X"20",
     X"aa", X"e7", X"a9", X"70", X"a0", X"f0", X"20", X"a7",
     X"e7", X"a5", X"a2", X"48", X"10", X"0d", X"20", X"a0",
     X"e7", X"a5", X"a2", X"30", X"09", X"a5", X"16", X"49",
     X"ff", X"85", X"16", X"20", X"d0", X"ee", X"a9", X"70",
     X"a0", X"f0", X"20", X"be", X"e7", X"68", X"10", X"03",
     X"20", X"d0", X"ee", X"a9", X"75", X"a0", X"f0", X"4c",
     X"5c", X"ef", X"20", X"21", X"eb", X"a9", X"00", X"85",
     X"16", X"20", X"f1", X"ef", X"a2", X"8a", X"a0", X"00",
     X"20", X"e7", X"ef", X"a9", X"93", X"a0", X"00", X"20",
     X"f9", X"ea", X"a9", X"00", X"85", X"a2", X"a5", X"16",
     X"20", X"62", X"f0", X"a9", X"8a", X"a0", X"00", X"4c",
     X"66", X"ea", X"48", X"4c", X"23", X"f0", X"81", X"49",
     X"0f", X"da", X"a2", X"83", X"49", X"0f", X"da", X"a2",
     X"7f", X"00", X"00", X"00", X"00", X"05", X"84", X"e6",
     X"1a", X"2d", X"1b", X"86", X"28", X"07", X"fb", X"f8",
     X"87", X"99", X"68", X"89", X"01", X"87", X"23", X"35",
     X"df", X"e1", X"86", X"a5", X"5d", X"e7", X"28", X"83",
     X"49", X"0f", X"da", X"a2", X"a6", X"d3", X"c1", X"c8",
     X"d4", X"c8", X"d5", X"c4", X"ce", X"ca", X"a5", X"a2",
     X"48", X"10", X"03", X"20", X"d0", X"ee", X"a5", X"9d",
     X"48", X"c9", X"81", X"90", X"07", X"a9", X"13", X"a0",
     X"e9", X"20", X"66", X"ea", X"a9", X"ce", X"a0", X"f0",
     X"20", X"5c", X"ef", X"68", X"c9", X"81", X"90", X"07",
     X"a9", X"66", X"a0", X"f0", X"20", X"a7", X"e7", X"68",
     X"10", X"03", X"4c", X"d0", X"ee", X"60", X"0b", X"76",
     X"b3", X"83", X"bd", X"d3", X"79", X"1e", X"f4", X"a6",
     X"f5", X"7b", X"83", X"fc", X"b0", X"10", X"7c", X"0c",
     X"1f", X"67", X"ca", X"7c", X"de", X"53", X"cb", X"c1",
     X"7d", X"14", X"64", X"70", X"4c", X"7d", X"b7", X"ea",
     X"51", X"7a", X"7d", X"63", X"30", X"88", X"7e", X"7e",
     X"92", X"44", X"99", X"3a", X"7e", X"4c", X"cc", X"91",
     X"c7", X"7f", X"aa", X"aa", X"aa", X"13", X"81", X"00",
     X"00", X"00", X"00", X"e6", X"b8", X"d0", X"02", X"e6",
     X"b9", X"ad", X"60", X"ea", X"c9", X"3a", X"b0", X"0a",
     X"c9", X"20", X"f0", X"ef", X"38", X"e9", X"30", X"38",
     X"e9", X"d0", X"60", X"80", X"4f", X"c7", X"52", X"58",
     X"a2", X"ff", X"86", X"76", X"a2", X"fb", X"9a", X"a9",
     X"28", X"a0", X"f1", X"85", X"01", X"84", X"02", X"85",
     X"04", X"84", X"05", X"20", X"73", X"f2", X"a9", X"4c",
     X"85", X"00", X"85", X"03", X"85", X"90", X"85", X"0a",
     X"a9", X"99", X"a0", X"e1", X"85", X"0b", X"84", X"0c",
     X"a2", X"1c", X"bd", X"0a", X"f1", X"95", X"b0", X"86",
     X"f1", X"ca", X"d0", X"f6", X"86", X"f2", X"8a", X"85",
     X"a4", X"85", X"54", X"48", X"a9", X"03", X"85", X"8f",
     X"20", X"fb", X"da", X"a9", X"01", X"8d", X"fd", X"01",
     X"8d", X"fc", X"01", X"a2", X"55", X"86", X"52", X"a9",
     X"00", X"a0", X"08", X"85", X"50", X"84", X"51", X"a0",
     X"00", X"e6", X"51", X"b1", X"50", X"49", X"ff", X"91",
     X"50", X"d1", X"50", X"d0", X"08", X"49", X"ff", X"91",
     X"50", X"d1", X"50", X"f0", X"ec", X"a4", X"50", X"a5",
     X"51", X"29", X"f0", X"84", X"73", X"85", X"74", X"84",
     X"6f", X"85", X"70", X"a2", X"00", X"a0", X"08", X"86",
     X"67", X"84", X"68", X"a0", X"00", X"84", X"d6", X"98",
     X"91", X"67", X"e6", X"67", X"d0", X"02", X"e6", X"68",
     X"a5", X"67", X"a4", X"68", X"20", X"e3", X"d3", X"20",
     X"4b", X"d6", X"a9", X"3a", X"a0", X"db", X"85", X"04",
     X"84", X"05", X"a9", X"3c", X"a0", X"d4", X"85", X"01",
     X"84", X"02", X"6c", X"01", X"00", X"20", X"67", X"dd",
     X"20", X"52", X"e7", X"6c", X"50", X"00", X"20", X"f8",
     X"e6", X"8a", X"4c", X"8b", X"fe", X"20", X"f8", X"e6",
     X"8a", X"4c", X"95", X"fe", X"20", X"f8", X"e6", X"e0",
     X"30", X"b0", X"13", X"86", X"f0", X"a9", X"2c", X"20",
     X"c0", X"de", X"20", X"f8", X"e6", X"e0", X"30", X"b0",
     X"05", X"86", X"2c", X"86", X"2d", X"60", X"4c", X"99",
     X"e1", X"20", X"ec", X"f1", X"e4", X"f0", X"b0", X"08",
     X"a5", X"f0", X"85", X"2c", X"85", X"2d", X"86", X"f0",
     X"a9", X"c5", X"20", X"c0", X"de", X"20", X"f8", X"e6",
     X"e0", X"30", X"b0", X"e2", X"60", X"20", X"ec", X"f1",
     X"8a", X"a4", X"f0", X"c0", X"28", X"b0", X"d7", X"4c",
     X"00", X"f8", X"20", X"09", X"f2", X"8a", X"a4", X"2c",
     X"c0", X"28", X"b0", X"ca", X"a4", X"f0", X"4c", X"19",
     X"f8", X"20", X"09", X"f2", X"8a", X"a8", X"c0", X"28",
     X"b0", X"bc", X"a5", X"f0", X"4c", X"28", X"f8", X"20",
     X"f8", X"e6", X"8a", X"4c", X"64", X"f8", X"20", X"f8",
     X"e6", X"ca", X"8a", X"c9", X"18", X"b0", X"a7", X"4c",
     X"5b", X"fb", X"20", X"f8", X"e6", X"8a", X"49", X"ff",
     X"aa", X"e8", X"86", X"f1", X"60", X"38", X"90", X"18",
     X"66", X"f2", X"60", X"a9", X"ff", X"d0", X"02", X"a9",
     X"3f", X"a2", X"00", X"85", X"32", X"86", X"f3", X"60",
     X"a9", X"7f", X"a2", X"40", X"d0", X"f5", X"20", X"67",
     X"dd", X"20", X"52", X"e7", X"a5", X"50", X"c5", X"6d",
     X"a5", X"51", X"e5", X"6e", X"b0", X"03", X"4c", X"10",
     X"d4", X"a5", X"50", X"85", X"73", X"85", X"6f", X"a5",
     X"51", X"85", X"74", X"85", X"70", X"60", X"20", X"67",
     X"dd", X"20", X"52", X"e7", X"a5", X"50", X"c5", X"73",
     X"a5", X"51", X"e5", X"74", X"b0", X"e0", X"a5", X"50",
     X"c5", X"69", X"a5", X"51", X"e5", X"6a", X"90", X"d6",
     X"a5", X"50", X"85", X"69", X"a5", X"51", X"85", X"6a",
     X"4c", X"6c", X"d6", X"a9", X"ab", X"20", X"c0", X"de",
     X"a5", X"b8", X"85", X"f4", X"a5", X"b9", X"85", X"f5",
     X"38", X"66", X"d8", X"a5", X"75", X"85", X"f6", X"a5",
     X"76", X"85", X"f7", X"20", X"a6", X"d9", X"4c", X"98",
     X"d9", X"86", X"de", X"a6", X"f8", X"86", X"df", X"a5",
     X"75", X"85", X"da", X"a5", X"76", X"85", X"db", X"a5",
     X"79", X"85", X"dc", X"a5", X"7a", X"85", X"dd", X"a5",
     X"f4", X"85", X"b8", X"a5", X"f5", X"85", X"b9", X"a5",
     X"f6", X"85", X"75", X"a5", X"f7", X"85", X"76", X"20",
     X"b7", X"00", X"20", X"3e", X"d9", X"4c", X"d2", X"d7",
     X"a5", X"da", X"85", X"75", X"a5", X"db", X"85", X"76",
     X"a5", X"dc", X"85", X"b8", X"a5", X"dd", X"85", X"b9",
     X"a6", X"df", X"9a", X"4c", X"d2", X"d7", X"4c", X"c9",
     X"de", X"b0", X"fb", X"a6", X"af", X"86", X"69", X"a6",
     X"b0", X"86", X"6a", X"20", X"0c", X"da", X"20", X"1a",
     X"d6", X"a5", X"9b", X"85", X"60", X"a5", X"9c", X"85",
     X"61", X"a9", X"2c", X"20", X"c0", X"de", X"20", X"0c",
     X"da", X"e6", X"50", X"d0", X"02", X"e6", X"51", X"20",
     X"1a", X"d6", X"a5", X"9b", X"c5", X"60", X"a5", X"9c",
     X"e5", X"61", X"b0", X"01", X"60", X"a0", X"00", X"b1",
     X"9b", X"91", X"60", X"e6", X"9b", X"d0", X"02", X"e6",
     X"9c", X"e6", X"60", X"d0", X"02", X"e6", X"61", X"a5",
     X"69", X"c5", X"9b", X"a5", X"6a", X"e5", X"9c", X"b0",
     X"e6", X"a6", X"61", X"a4", X"60", X"d0", X"01", X"ca",
     X"88", X"86", X"6a", X"84", X"69", X"4c", X"f2", X"d4",
     X"ad", X"56", X"c0", X"ad", X"53", X"c0", X"4c", X"40",
     X"fb", X"ad", X"54", X"c0", X"4c", X"39", X"fb", X"20",
     X"d9", X"f7", X"a0", X"03", X"b1", X"9b", X"aa", X"88",
     X"b1", X"9b", X"e9", X"01", X"b0", X"01", X"ca", X"85",
     X"50", X"86", X"51", X"20", X"cd", X"fe", X"20", X"bc",
     X"f7", X"4c", X"cd", X"fe", X"20", X"d9", X"f7", X"20",
     X"fd", X"fe", X"a0", X"02", X"b1", X"9b", X"c5", X"50",
     X"c8", X"b1", X"9b", X"e5", X"51", X"b0", X"03", X"4c",
     X"10", X"d4", X"20", X"bc", X"f7", X"4c", X"fd", X"fe",
     X"2c", X"55", X"c0", X"2c", X"52", X"c0", X"a9", X"40",
     X"d0", X"08", X"a9", X"20", X"2c", X"54", X"c0", X"2c",
     X"53", X"c0", X"85", X"e6", X"ad", X"57", X"c0", X"ad",
     X"50", X"c0", X"a9", X"00", X"85", X"1c", X"a5", X"e6",
     X"85", X"1b", X"a0", X"00", X"84", X"1a", X"a5", X"1c",
     X"91", X"1a", X"20", X"7e", X"f4", X"c8", X"d0", X"f6",
     X"e6", X"1b", X"a5", X"1b", X"29", X"1f", X"d0", X"ee",
     X"60", X"85", X"e2", X"86", X"e0", X"84", X"e1", X"48",
     X"29", X"c0", X"85", X"26", X"4a", X"4a", X"05", X"26",
     X"85", X"26", X"68", X"85", X"27", X"0a", X"0a", X"0a",
     X"26", X"27", X"0a", X"26", X"27", X"0a", X"66", X"26",
     X"a5", X"27", X"29", X"1f", X"05", X"e6", X"85", X"27",
     X"8a", X"c0", X"00", X"f0", X"05", X"a0", X"23", X"69",
     X"04", X"c8", X"e9", X"07", X"b0", X"fb", X"84", X"e5",
     X"aa", X"bd", X"b9", X"f4", X"85", X"30", X"98", X"4a",
     X"a5", X"e4", X"85", X"1c", X"b0", X"28", X"60", X"20",
     X"11", X"f4", X"a5", X"1c", X"51", X"26", X"25", X"30",
     X"51", X"26", X"91", X"26", X"60", X"10", X"23", X"a5",
     X"30", X"4a", X"b0", X"05", X"49", X"c0", X"85", X"30",
     X"60", X"88", X"10", X"02", X"a0", X"27", X"a9", X"c0",
     X"85", X"30", X"84", X"e5", X"a5", X"1c", X"0a", X"c9",
     X"c0", X"10", X"06", X"a5", X"1c", X"49", X"7f", X"85",
     X"1c", X"60", X"a5", X"30", X"0a", X"49", X"80", X"30",
     X"dd", X"a9", X"81", X"c8", X"c0", X"28", X"90", X"e0",
     X"a0", X"00", X"b0", X"dc", X"18", X"a5", X"d1", X"29",
     X"04", X"f0", X"25", X"a9", X"7f", X"25", X"30", X"31",
     X"26", X"d0", X"19", X"e6", X"ea", X"a9", X"7f", X"25",
     X"30", X"10", X"11", X"18", X"a5", X"d1", X"29", X"04",
     X"f0", X"0e", X"b1", X"26", X"45", X"1c", X"25", X"30",
     X"d0", X"02", X"e6", X"ea", X"51", X"26", X"91", X"26",
     X"a5", X"d1", X"65", X"d3", X"29", X"03", X"c9", X"02",
     X"6a", X"b0", X"92", X"30", X"30", X"18", X"a5", X"27",
     X"2c", X"b9", X"f5", X"d0", X"22", X"06", X"26", X"b0",
     X"1a", X"2c", X"cd", X"f4", X"f0", X"05", X"69", X"1f",
     X"38", X"b0", X"12", X"69", X"23", X"48", X"a5", X"26",
     X"69", X"b0", X"b0", X"02", X"69", X"f0", X"85", X"26",
     X"68", X"b0", X"02", X"69", X"1f", X"66", X"26", X"69",
     X"fc", X"85", X"27", X"60", X"18", X"a5", X"27", X"69",
     X"04", X"2c", X"b9", X"f5", X"d0", X"f3", X"06", X"26",
     X"90", X"18", X"69", X"e0", X"18", X"2c", X"08", X"f5",
     X"f0", X"12", X"a5", X"26", X"69", X"50", X"49", X"f0",
     X"f0", X"02", X"49", X"f0", X"85", X"26", X"a5", X"e6",
     X"90", X"02", X"69", X"e0", X"66", X"26", X"90", X"d1",
     X"48", X"a9", X"00", X"85", X"e0", X"85", X"e1", X"85",
     X"e2", X"68", X"48", X"38", X"e5", X"e0", X"48", X"8a",
     X"e5", X"e1", X"85", X"d3", X"b0", X"0a", X"68", X"49",
     X"ff", X"69", X"01", X"48", X"a9", X"00", X"e5", X"d3",
     X"85", X"d1", X"85", X"d5", X"68", X"85", X"d0", X"85",
     X"d4", X"68", X"85", X"e0", X"86", X"e1", X"98", X"18",
     X"e5", X"e2", X"90", X"04", X"49", X"ff", X"69", X"fe",
     X"85", X"d2", X"84", X"e2", X"66", X"d3", X"38", X"e5",
     X"d0", X"aa", X"a9", X"ff", X"e5", X"d1", X"85", X"1d",
     X"a4", X"e5", X"b0", X"05", X"0a", X"20", X"65", X"f4",
     X"38", X"a5", X"d4", X"65", X"d2", X"85", X"d4", X"a5",
     X"d5", X"e9", X"00", X"85", X"d5", X"b1", X"26", X"45",
     X"1c", X"25", X"30", X"51", X"26", X"91", X"26", X"e8",
     X"d0", X"04", X"e6", X"1d", X"f0", X"62", X"a5", X"d3",
     X"b0", X"da", X"20", X"d3", X"f4", X"18", X"a5", X"d4",
     X"65", X"d0", X"85", X"d4", X"a5", X"d5", X"65", X"d1",
     X"50", X"d9", X"81", X"82", X"84", X"88", X"90", X"a0",
     X"c0", X"1c", X"ff", X"fe", X"fa", X"f4", X"ec", X"e1",
     X"d4", X"c5", X"b4", X"a1", X"8d", X"78", X"61", X"49",
     X"31", X"18", X"ff", X"a5", X"26", X"0a", X"a5", X"27",
     X"29", X"03", X"2a", X"05", X"26", X"0a", X"0a", X"0a",
     X"85", X"e2", X"a5", X"27", X"4a", X"4a", X"29", X"07",
     X"05", X"e2", X"85", X"e2", X"a5", X"e5", X"0a", X"65",
     X"e5", X"0a", X"aa", X"ca", X"a5", X"30", X"29", X"7f",
     X"e8", X"4a", X"d0", X"fc", X"85", X"e1", X"8a", X"18",
     X"65", X"e5", X"90", X"02", X"e6", X"e1", X"85", X"e0",
     X"60", X"86", X"1a", X"84", X"1b", X"aa", X"4a", X"4a",
     X"4a", X"4a", X"85", X"d3", X"8a", X"29", X"0f", X"aa",
     X"bc", X"ba", X"f5", X"84", X"d0", X"49", X"0f", X"aa",
     X"bc", X"bb", X"f5", X"c8", X"84", X"d2", X"a4", X"e5",
     X"a2", X"00", X"86", X"ea", X"a1", X"1a", X"85", X"d1",
     X"a2", X"80", X"86", X"d4", X"86", X"d5", X"a6", X"e7",
     X"a5", X"d4", X"38", X"65", X"d0", X"85", X"d4", X"90",
     X"04", X"20", X"b3", X"f4", X"18", X"a5", X"d5", X"65",
     X"d2", X"85", X"d5", X"90", X"03", X"20", X"b4", X"f4",
     X"ca", X"d0", X"e5", X"a5", X"d1", X"4a", X"4a", X"4a",
     X"d0", X"d4", X"e6", X"1a", X"d0", X"02", X"e6", X"1b",
     X"a1", X"1a", X"d0", X"ca", X"60", X"86", X"1a", X"84",
     X"1b", X"aa", X"4a", X"4a", X"4a", X"4a", X"85", X"d3",
     X"8a", X"29", X"0f", X"aa", X"bc", X"ba", X"f5", X"84",
     X"d0", X"49", X"0f", X"aa", X"bc", X"bb", X"f5", X"c8",
     X"84", X"d2", X"a4", X"e5", X"a2", X"00", X"86", X"ea",
     X"a1", X"1a", X"85", X"d1", X"a2", X"80", X"86", X"d4",
     X"86", X"d5", X"a6", X"e7", X"a5", X"d4", X"38", X"65",
     X"d0", X"85", X"d4", X"90", X"04", X"20", X"9c", X"f4",
     X"18", X"a5", X"d5", X"65", X"d2", X"85", X"d5", X"90",
     X"03", X"20", X"9d", X"f4", X"ca", X"d0", X"e5", X"a5",
     X"d1", X"4a", X"4a", X"4a", X"d0", X"d4", X"e6", X"1a",
     X"d0", X"02", X"e6", X"1b", X"a1", X"1a", X"d0", X"ca",
     X"60", X"20", X"67", X"dd", X"20", X"52", X"e7", X"a4",
     X"51", X"a6", X"50", X"c0", X"01", X"90", X"06", X"d0",
     X"1d", X"e0", X"18", X"b0", X"19", X"8a", X"48", X"98",
     X"48", X"a9", X"2c", X"20", X"c0", X"de", X"20", X"f8",
     X"e6", X"e0", X"c0", X"b0", X"09", X"86", X"9d", X"68",
     X"a8", X"68", X"aa", X"a5", X"9d", X"60", X"4c", X"06",
     X"f2", X"20", X"f8", X"e6", X"e0", X"08", X"b0", X"f6",
     X"bd", X"f6", X"f6", X"85", X"e4", X"60", X"00", X"2a",
     X"55", X"7f", X"80", X"aa", X"d5", X"ff", X"c9", X"c1",
     X"f0", X"0d", X"20", X"b9", X"f6", X"20", X"57", X"f4",
     X"20", X"b7", X"00", X"c9", X"c1", X"d0", X"e6", X"20",
     X"c0", X"de", X"20", X"b9", X"f6", X"84", X"9d", X"a8",
     X"8a", X"a6", X"9d", X"20", X"3a", X"f5", X"4c", X"08",
     X"f7", X"20", X"f8", X"e6", X"86", X"f9", X"60", X"20",
     X"f8", X"e6", X"86", X"e7", X"60", X"20", X"f8", X"e6",
     X"a5", X"e8", X"85", X"1a", X"a5", X"e9", X"85", X"1b",
     X"8a", X"a2", X"00", X"c1", X"1a", X"f0", X"02", X"b0",
     X"a5", X"0a", X"90", X"03", X"e6", X"1b", X"18", X"a8",
     X"b1", X"1a", X"65", X"1a", X"aa", X"c8", X"b1", X"1a",
     X"65", X"e9", X"85", X"1b", X"86", X"1a", X"20", X"b7",
     X"00", X"c9", X"c5", X"d0", X"09", X"20", X"c0", X"de",
     X"20", X"b9", X"f6", X"20", X"11", X"f4", X"a5", X"f9",
     X"60", X"20", X"2d", X"f7", X"4c", X"05", X"f6", X"20",
     X"2d", X"f7", X"4c", X"61", X"f6", X"a9", X"00", X"85",
     X"3d", X"85", X"3f", X"a0", X"50", X"84", X"3c", X"c8",
     X"84", X"3e", X"20", X"fd", X"fe", X"18", X"a5", X"73",
     X"aa", X"ca", X"86", X"3e", X"e5", X"50", X"48", X"a5",
     X"74", X"a8", X"e8", X"d0", X"01", X"88", X"84", X"3f",
     X"e5", X"51", X"c5", X"6e", X"90", X"02", X"d0", X"03",
     X"4c", X"10", X"d4", X"85", X"74", X"85", X"70", X"85",
     X"3d", X"85", X"e9", X"68", X"85", X"e8", X"85", X"73",
     X"85", X"6f", X"85", X"3c", X"20", X"fa", X"fc", X"a9",
     X"03", X"4c", X"02", X"ff", X"18", X"a5", X"9b", X"65",
     X"50", X"85", X"3e", X"a5", X"9c", X"65", X"51", X"85",
     X"3f", X"a0", X"04", X"b1", X"9b", X"20", X"ef", X"e0",
     X"a5", X"94", X"85", X"3c", X"a5", X"95", X"85", X"3d",
     X"60", X"a9", X"40", X"85", X"14", X"20", X"e3", X"df",
     X"a9", X"00", X"85", X"14", X"4c", X"f0", X"d8", X"20",
     X"f8", X"e6", X"ca", X"8a", X"c9", X"28", X"90", X"0a",
     X"e9", X"28", X"48", X"20", X"fb", X"da", X"68", X"4c",
     X"ec", X"f7", X"85", X"24", X"60", X"cb", X"d2", X"d7",
     X"4a", X"08", X"20", X"47", X"f8", X"28", X"a9", X"0f",
     X"90", X"02", X"69", X"e0", X"85", X"2e", X"b1", X"26",
     X"45", X"30", X"25", X"2e", X"51", X"26", X"91", X"26",
     X"60", X"20", X"00", X"f8", X"c4", X"2c", X"b0", X"11",
     X"c8", X"20", X"0e", X"f8", X"90", X"f6", X"69", X"01",
     X"48", X"20", X"00", X"f8", X"68", X"c5", X"2d", X"90",
     X"f5", X"60", X"a0", X"2f", X"d0", X"02", X"a0", X"27",
     X"84", X"2d", X"a0", X"27", X"a9", X"00", X"85", X"30",
     X"20", X"28", X"f8", X"88", X"10", X"f6", X"60", X"48",
     X"4a", X"29", X"03", X"09", X"04", X"85", X"27", X"68",
     X"29", X"18", X"90", X"02", X"69", X"7f", X"85", X"26",
     X"0a", X"0a", X"05", X"26", X"85", X"26", X"60", X"a5",
     X"30", X"18", X"69", X"03", X"29", X"0f", X"85", X"30",
     X"0a", X"0a", X"0a", X"0a", X"05", X"30", X"85", X"30",
     X"60", X"4a", X"08", X"20", X"47", X"f8", X"b1", X"26",
     X"28", X"90", X"04", X"4a", X"4a", X"4a", X"4a", X"29",
     X"0f", X"60", X"a6", X"3a", X"a4", X"3b", X"20", X"96",
     X"fd", X"20", X"48", X"f9", X"a1", X"3a", X"a8", X"4a",
     X"90", X"09", X"6a", X"b0", X"10", X"c9", X"a2", X"f0",
     X"0c", X"29", X"87", X"4a", X"aa", X"bd", X"62", X"f9",
     X"20", X"79", X"f8", X"d0", X"04", X"a0", X"80", X"a9",
     X"00", X"aa", X"bd", X"a6", X"f9", X"85", X"2e", X"29",
     X"03", X"85", X"2f", X"98", X"29", X"8f", X"aa", X"98",
     X"a0", X"03", X"e0", X"8a", X"f0", X"0b", X"4a", X"90",
     X"08", X"4a", X"4a", X"09", X"20", X"88", X"d0", X"fa",
     X"c8", X"88", X"d0", X"f2", X"60", X"ff", X"ff", X"ff",
     X"20", X"82", X"f8", X"48", X"b1", X"3a", X"20", X"da",
     X"fd", X"a2", X"01", X"20", X"4a", X"f9", X"c4", X"2f",
     X"c8", X"90", X"f1", X"a2", X"03", X"c0", X"04", X"90",
     X"f2", X"68", X"a8", X"b9", X"c0", X"f9", X"85", X"2c",
     X"b9", X"00", X"fa", X"85", X"2d", X"a9", X"00", X"a0",
     X"05", X"06", X"2d", X"26", X"2c", X"2a", X"88", X"d0",
     X"f8", X"69", X"bf", X"20", X"ed", X"fd", X"ca", X"d0",
     X"ec", X"20", X"48", X"f9", X"a4", X"2f", X"a2", X"06",
     X"e0", X"03", X"f0", X"1c", X"06", X"2e", X"90", X"0e",
     X"bd", X"b3", X"f9", X"20", X"ed", X"fd", X"bd", X"b9",
     X"f9", X"f0", X"03", X"20", X"ed", X"fd", X"ca", X"d0",
     X"e7", X"60", X"88", X"30", X"e7", X"20", X"da", X"fd",
     X"a5", X"2e", X"c9", X"e8", X"b1", X"3a", X"90", X"f2",
     X"20", X"56", X"f9", X"aa", X"e8", X"d0", X"01", X"c8",
     X"98", X"20", X"da", X"fd", X"8a", X"4c", X"da", X"fd",
     X"a2", X"03", X"a9", X"a0", X"20", X"ed", X"fd", X"ca",
     X"d0", X"f8", X"60", X"38", X"a5", X"2f", X"a4", X"3b",
     X"aa", X"10", X"01", X"88", X"65", X"3a", X"90", X"01",
     X"c8", X"60", X"04", X"20", X"54", X"30", X"0d", X"80",
     X"04", X"90", X"03", X"22", X"54", X"33", X"0d", X"80",
     X"04", X"90", X"04", X"20", X"54", X"33", X"0d", X"80",
     X"04", X"90", X"04", X"20", X"54", X"3b", X"0d", X"80",
     X"04", X"90", X"00", X"22", X"44", X"33", X"0d", X"c8",
     X"44", X"00", X"11", X"22", X"44", X"33", X"0d", X"c8",
     X"44", X"a9", X"01", X"22", X"44", X"33", X"0d", X"80",
     X"04", X"90", X"01", X"22", X"44", X"33", X"0d", X"80",
     X"04", X"90", X"26", X"31", X"87", X"9a", X"00", X"21",
     X"81", X"82", X"00", X"00", X"59", X"4d", X"91", X"92",
     X"86", X"4a", X"85", X"9d", X"ac", X"a9", X"ac", X"a3",
     X"a8", X"a4", X"d9", X"00", X"d8", X"a4", X"a4", X"00",
     X"1c", X"8a", X"1c", X"23", X"5d", X"8b", X"1b", X"a1",
     X"9d", X"8a", X"1d", X"23", X"9d", X"8b", X"1d", X"a1",
     X"00", X"29", X"19", X"ae", X"69", X"a8", X"19", X"23",
     X"24", X"53", X"1b", X"23", X"24", X"53", X"19", X"a1",
     X"00", X"1a", X"5b", X"5b", X"a5", X"69", X"24", X"24",
     X"ae", X"ae", X"a8", X"ad", X"29", X"00", X"7c", X"00",
     X"15", X"9c", X"6d", X"9c", X"a5", X"69", X"29", X"53",
     X"84", X"13", X"34", X"11", X"a5", X"69", X"23", X"a0",
     X"d8", X"62", X"5a", X"48", X"26", X"62", X"94", X"88",
     X"54", X"44", X"c8", X"54", X"68", X"44", X"e8", X"94",
     X"00", X"b4", X"08", X"84", X"74", X"b4", X"28", X"6e",
     X"74", X"f4", X"cc", X"4a", X"72", X"f2", X"a4", X"8a",
     X"00", X"aa", X"a2", X"a2", X"74", X"74", X"74", X"72",
     X"44", X"68", X"b2", X"32", X"b2", X"00", X"22", X"00",
     X"1a", X"1a", X"26", X"26", X"72", X"72", X"88", X"c8",
     X"c4", X"ca", X"26", X"48", X"44", X"44", X"a2", X"c8",
     X"85", X"45", X"68", X"48", X"0a", X"0a", X"0a", X"30",
     X"03", X"6c", X"fe", X"03", X"28", X"20", X"4c", X"ff",
     X"68", X"85", X"3a", X"68", X"85", X"3b", X"6c", X"f0",
     X"03", X"20", X"82", X"f8", X"20", X"da", X"fa", X"4c",
     X"65", X"ff", X"d8", X"20", X"84", X"fe", X"20", X"2f",
     X"fb", X"20", X"93", X"fe", X"20", X"89", X"fe", X"ad",
     X"58", X"c0", X"ad", X"5a", X"c0", X"ad", X"5d", X"c0",
     X"ad", X"5f", X"c0", X"ad", X"ff", X"cf", X"2c", X"10",
     X"c0", X"d8", X"20", X"3a", X"ff", X"ad", X"f3", X"03",
     X"49", X"a5", X"cd", X"f4", X"03", X"d0", X"17", X"ad",
     X"f2", X"03", X"d0", X"0f", X"a9", X"e0", X"cd", X"f3",
     X"03", X"d0", X"08", X"a0", X"03", X"8c", X"f2", X"03",
     X"4c", X"00", X"e0", X"6c", X"f2", X"03", X"20", X"60",
     X"fb", X"a2", X"05", X"bd", X"fc", X"fa", X"9d", X"ef",
     X"03", X"ca", X"d0", X"f7", X"a9", X"c8", X"86", X"00",
     X"85", X"01", X"a0", X"07", X"c6", X"01", X"a5", X"01",
     X"c9", X"c0", X"f0", X"d7", X"8d", X"f8", X"07", X"b1",
     X"00", X"d9", X"01", X"fb", X"d0", X"ec", X"88", X"88",
     X"10", X"f5", X"6c", X"00", X"00", X"ea", X"ea", X"20",
     X"8e", X"fd", X"a9", X"45", X"85", X"40", X"a9", X"00",
     X"85", X"41", X"a2", X"fb", X"a9", X"a0", X"20", X"ed",
     X"fd", X"bd", X"1e", X"fa", X"20", X"ed", X"fd", X"a9",
     X"bd", X"20", X"ed", X"fd", X"b5", X"4a", X"20", X"da",
     X"fd", X"e8", X"30", X"e8", X"60", X"59", X"fa", X"00",
     X"e0", X"45", X"20", X"ff", X"00", X"ff", X"03", X"ff",
     X"3c", X"c1", X"d0", X"d0", X"cc", X"c5", X"a0", X"dd",
     X"db", X"c4", X"c2", X"c1", X"ff", X"c3", X"ff", X"ff",
     X"ff", X"c1", X"d8", X"d9", X"d0", X"d3", X"ad", X"70",
     X"c0", X"a0", X"00", X"ea", X"ea", X"bd", X"64", X"c0",
     X"10", X"04", X"c8", X"d0", X"f8", X"88", X"60", X"a9",
     X"00", X"85", X"48", X"ad", X"56", X"c0", X"ad", X"54",
     X"c0", X"ad", X"51", X"c0", X"a9", X"00", X"f0", X"0b",
     X"ad", X"50", X"c0", X"ad", X"53", X"c0", X"20", X"36",
     X"f8", X"a9", X"14", X"85", X"22", X"a9", X"00", X"85",
     X"20", X"a9", X"28", X"85", X"21", X"a9", X"18", X"85",
     X"23", X"a9", X"17", X"85", X"25", X"4c", X"22", X"fc",
     X"20", X"58", X"fc", X"a0", X"08", X"b9", X"08", X"fb",
     X"99", X"0e", X"04", X"88", X"d0", X"f7", X"60", X"ad",
     X"f3", X"03", X"49", X"a5", X"8d", X"f4", X"03", X"60",
     X"c9", X"8d", X"d0", X"18", X"ac", X"00", X"c0", X"10",
     X"13", X"c0", X"93", X"d0", X"0f", X"2c", X"10", X"c0",
     X"ac", X"00", X"c0", X"10", X"fb", X"c0", X"83", X"f0",
     X"03", X"2c", X"10", X"c0", X"4c", X"fd", X"fb", X"38",
     X"4c", X"2c", X"fc", X"a8", X"b9", X"48", X"fa", X"20",
     X"97", X"fb", X"20", X"0c", X"fd", X"c9", X"ce", X"b0",
     X"ee", X"c9", X"c9", X"90", X"ea", X"c9", X"cc", X"f0",
     X"e6", X"d0", X"e8", X"ea", X"ea", X"ea", X"ea", X"ea",
     X"ea", X"ea", X"ea", X"ea", X"ea", X"ea", X"ea", X"ea",
     X"ea", X"48", X"4a", X"29", X"03", X"09", X"04", X"85",
     X"29", X"68", X"29", X"18", X"90", X"02", X"69", X"7f",
     X"85", X"28", X"0a", X"0a", X"05", X"28", X"85", X"28",
     X"60", X"c9", X"87", X"d0", X"12", X"a9", X"40", X"20",
     X"a8", X"fc", X"a0", X"c0", X"a9", X"0c", X"20", X"a8",
     X"fc", X"ad", X"30", X"c0", X"88", X"d0", X"f5", X"60",
     X"a4", X"24", X"91", X"28", X"e6", X"24", X"a5", X"24",
     X"c5", X"21", X"b0", X"66", X"60", X"c9", X"a0", X"b0",
     X"ef", X"a8", X"10", X"ec", X"c9", X"8d", X"f0", X"5a",
     X"c9", X"8a", X"f0", X"5a", X"c9", X"88", X"d0", X"c9",
     X"c6", X"24", X"10", X"e8", X"a5", X"21", X"85", X"24",
     X"c6", X"24", X"a5", X"22", X"c5", X"25", X"b0", X"0b",
     X"c6", X"25", X"a5", X"25", X"20", X"c1", X"fb", X"65",
     X"20", X"85", X"28", X"60", X"49", X"c0", X"f0", X"28",
     X"69", X"fd", X"90", X"c0", X"f0", X"da", X"69", X"fd",
     X"90", X"2c", X"f0", X"de", X"69", X"fd", X"90", X"5c",
     X"d0", X"e9", X"a4", X"24", X"a5", X"25", X"48", X"20",
     X"24", X"fc", X"20", X"9e", X"fc", X"a0", X"00", X"68",
     X"69", X"00", X"c5", X"23", X"90", X"f0", X"b0", X"ca",
     X"a5", X"22", X"85", X"25", X"a0", X"00", X"84", X"24",
     X"f0", X"e4", X"a9", X"00", X"85", X"24", X"e6", X"25",
     X"a5", X"25", X"c5", X"23", X"90", X"b6", X"c6", X"25",
     X"a5", X"22", X"48", X"20", X"24", X"fc", X"a5", X"28",
     X"85", X"2a", X"a5", X"29", X"85", X"2b", X"a4", X"21",
     X"88", X"68", X"69", X"01", X"c5", X"23", X"b0", X"0d",
     X"48", X"20", X"24", X"fc", X"b1", X"28", X"91", X"2a",
     X"88", X"10", X"f9", X"30", X"e1", X"a0", X"00", X"20",
     X"9e", X"fc", X"b0", X"86", X"a4", X"24", X"a9", X"a0",
     X"91", X"28", X"c8", X"c4", X"21", X"90", X"f9", X"60",
     X"38", X"48", X"e9", X"01", X"d0", X"fc", X"68", X"e9",
     X"01", X"d0", X"f6", X"60", X"e6", X"42", X"d0", X"02",
     X"e6", X"43", X"a5", X"3c", X"c5", X"3e", X"a5", X"3d",
     X"e5", X"3f", X"e6", X"3c", X"d0", X"02", X"e6", X"3d",
     X"60", X"a0", X"4b", X"20", X"db", X"fc", X"d0", X"f9",
     X"69", X"fe", X"b0", X"f5", X"a0", X"21", X"20", X"db",
     X"fc", X"c8", X"c8", X"88", X"d0", X"fd", X"90", X"05",
     X"a0", X"32", X"88", X"d0", X"fd", X"ac", X"20", X"c0",
     X"a0", X"2c", X"ca", X"60", X"a2", X"08", X"48", X"20",
     X"fa", X"fc", X"68", X"2a", X"a0", X"3a", X"ca", X"d0",
     X"f5", X"60", X"20", X"fd", X"fc", X"88", X"ad", X"60",
     X"c0", X"45", X"2f", X"10", X"f8", X"45", X"2f", X"85",
     X"2f", X"c0", X"80", X"60", X"a4", X"24", X"b1", X"28",
     X"48", X"29", X"3f", X"09", X"40", X"91", X"28", X"68",
     X"6c", X"38", X"00", X"e6", X"4e", X"d0", X"02", X"e6",
     X"4f", X"2c", X"00", X"c0", X"10", X"f5", X"91", X"28",
     X"ad", X"00", X"c0", X"2c", X"10", X"c0", X"60", X"20",
     X"0c", X"fd", X"20", X"a5", X"fb", X"20", X"0c", X"fd",
     X"c9", X"9b", X"f0", X"f3", X"60", X"a5", X"32", X"48",
     X"a9", X"ff", X"85", X"32", X"bd", X"00", X"02", X"20",
     X"ed", X"fd", X"68", X"85", X"32", X"bd", X"00", X"02",
     X"c9", X"88", X"f0", X"1d", X"c9", X"98", X"f0", X"0a",
     X"e0", X"f8", X"90", X"03", X"20", X"3a", X"ff", X"e8",
     X"d0", X"13", X"a9", X"dc", X"20", X"ed", X"fd", X"20",
     X"8e", X"fd", X"a5", X"33", X"20", X"ed", X"fd", X"a2",
     X"01", X"8a", X"f0", X"f3", X"ca", X"20", X"35", X"fd",
     X"c9", X"95", X"d0", X"02", X"b1", X"28", X"c9", X"e0",
     X"90", X"02", X"29", X"df", X"9d", X"00", X"02", X"c9",
     X"8d", X"d0", X"b2", X"20", X"9c", X"fc", X"a9", X"8d",
     X"d0", X"5b", X"a4", X"3d", X"a6", X"3c", X"20", X"8e",
     X"fd", X"20", X"40", X"f9", X"a0", X"00", X"a9", X"ad",
     X"4c", X"ed", X"fd", X"a5", X"3c", X"09", X"07", X"85",
     X"3e", X"a5", X"3d", X"85", X"3f", X"a5", X"3c", X"29",
     X"07", X"d0", X"03", X"20", X"92", X"fd", X"a9", X"a0",
     X"20", X"ed", X"fd", X"b1", X"3c", X"20", X"da", X"fd",
     X"20", X"ba", X"fc", X"90", X"e8", X"60", X"4a", X"90",
     X"ea", X"4a", X"4a", X"a5", X"3e", X"90", X"02", X"49",
     X"ff", X"65", X"3c", X"48", X"a9", X"bd", X"20", X"ed",
     X"fd", X"68", X"48", X"4a", X"4a", X"4a", X"4a", X"20",
     X"e5", X"fd", X"68", X"29", X"0f", X"09", X"b0", X"c9",
     X"ba", X"90", X"02", X"69", X"06", X"6c", X"36", X"00",
     X"c9", X"a0", X"90", X"02", X"25", X"32", X"84", X"35",
     X"48", X"20", X"78", X"fb", X"68", X"a4", X"35", X"60",
     X"c6", X"34", X"f0", X"9f", X"ca", X"d0", X"16", X"c9",
     X"ba", X"d0", X"bb", X"85", X"31", X"a5", X"3e", X"91",
     X"40", X"e6", X"40", X"d0", X"02", X"e6", X"41", X"60",
     X"a4", X"34", X"b9", X"ff", X"01", X"85", X"31", X"60",
     X"a2", X"01", X"b5", X"3e", X"95", X"42", X"95", X"44",
     X"ca", X"10", X"f7", X"60", X"b1", X"3c", X"91", X"42",
     X"20", X"b4", X"fc", X"90", X"f7", X"60", X"b1", X"3c",
     X"d1", X"42", X"f0", X"1c", X"20", X"92", X"fd", X"b1",
     X"3c", X"20", X"da", X"fd", X"a9", X"a0", X"20", X"ed",
     X"fd", X"a9", X"a8", X"20", X"ed", X"fd", X"b1", X"42",
     X"20", X"da", X"fd", X"a9", X"a9", X"20", X"ed", X"fd",
     X"20", X"b4", X"fc", X"90", X"d9", X"60", X"20", X"75",
     X"fe", X"a9", X"14", X"48", X"20", X"d0", X"f8", X"20",
     X"53", X"f9", X"85", X"3a", X"84", X"3b", X"68", X"38",
     X"e9", X"01", X"d0", X"ef", X"60", X"8a", X"f0", X"07",
     X"b5", X"3c", X"95", X"3a", X"ca", X"10", X"f9", X"60",
     X"a0", X"3f", X"d0", X"02", X"a0", X"ff", X"84", X"32",
     X"60", X"a9", X"00", X"85", X"3e", X"a2", X"38", X"a0",
     X"1b", X"d0", X"08", X"a9", X"00", X"85", X"3e", X"a2",
     X"36", X"a0", X"f0", X"a5", X"3e", X"29", X"0f", X"f0",
     X"06", X"09", X"c0", X"a0", X"00", X"f0", X"02", X"a9",
     X"fd", X"94", X"00", X"95", X"01", X"60", X"ea", X"ea",
     X"4c", X"00", X"e0", X"4c", X"03", X"e0", X"20", X"75",
     X"fe", X"20", X"3f", X"ff", X"6c", X"3a", X"00", X"4c",
     X"d7", X"fa", X"60", X"ea", X"60", X"ea", X"ea", X"ea",
     X"ea", X"ea", X"4c", X"f8", X"03", X"a9", X"40", X"20",
     X"c9", X"fc", X"a0", X"27", X"a2", X"00", X"41", X"3c",
     X"48", X"a1", X"3c", X"20", X"ed", X"fe", X"20", X"ba",
     X"fc", X"a0", X"1d", X"68", X"90", X"ee", X"a0", X"22",
     X"20", X"ed", X"fe", X"f0", X"4d", X"a2", X"10", X"0a",
     X"20", X"d6", X"fc", X"d0", X"fa", X"60", X"20", X"00",
     X"fe", X"68", X"68", X"d0", X"6c", X"20", X"fa", X"fc",
     X"a9", X"16", X"20", X"c9", X"fc", X"85", X"2e", X"20",
     X"fa", X"fc", X"a0", X"24", X"20", X"fd", X"fc", X"b0",
     X"f9", X"20", X"fd", X"fc", X"a0", X"3b", X"20", X"ec",
     X"fc", X"81", X"3c", X"45", X"2e", X"85", X"2e", X"20",
     X"ba", X"fc", X"a0", X"35", X"90", X"f0", X"20", X"ec",
     X"fc", X"c5", X"2e", X"f0", X"0d", X"a9", X"c5", X"20",
     X"ed", X"fd", X"a9", X"d2", X"20", X"ed", X"fd", X"20",
     X"ed", X"fd", X"a9", X"87", X"4c", X"ed", X"fd", X"a5",
     X"48", X"48", X"a5", X"45", X"a6", X"46", X"a4", X"47",
     X"28", X"60", X"85", X"45", X"86", X"46", X"84", X"47",
     X"08", X"68", X"85", X"48", X"ba", X"86", X"49", X"d8",
     X"60", X"20", X"84", X"fe", X"20", X"2f", X"fb", X"20",
     X"93", X"fe", X"20", X"89", X"fe", X"d8", X"20", X"3a",
     X"ff", X"a9", X"aa", X"85", X"33", X"20", X"67", X"fd",
     X"20", X"c7", X"ff", X"20", X"a7", X"ff", X"84", X"34",
     X"a0", X"17", X"88", X"30", X"e8", X"d9", X"cc", X"ff",
     X"d0", X"f8", X"20", X"be", X"ff", X"a4", X"34", X"4c",
     X"73", X"ff", X"a2", X"03", X"0a", X"0a", X"0a", X"0a",
     X"0a", X"26", X"3e", X"26", X"3f", X"ca", X"10", X"f8",
     X"a5", X"31", X"d0", X"06", X"b5", X"3f", X"95", X"3d",
     X"95", X"41", X"e8", X"f0", X"f3", X"d0", X"06", X"a2",
     X"00", X"86", X"3e", X"86", X"3f", X"b9", X"00", X"02",
     X"c8", X"49", X"b0", X"c9", X"0a", X"90", X"d3", X"69",
     X"88", X"c9", X"fa", X"b0", X"cd", X"60", X"a9", X"fe",
     X"48", X"b9", X"e3", X"ff", X"48", X"a5", X"31", X"a0",
     X"00", X"84", X"31", X"60", X"bc", X"b2", X"be", X"b2",
     X"ef", X"c4", X"b2", X"a9", X"bb", X"a6", X"a4", X"06",
     X"95", X"07", X"02", X"05", X"f0", X"00", X"eb", X"93",
     X"a7", X"c6", X"99", X"b2", X"c9", X"be", X"c1", X"35",
     X"8c", X"c4", X"96", X"af", X"17", X"17", X"2b", X"1f",
     X"83", X"7f", X"5d", X"cc", X"b5", X"fc", X"17", X"17",
     X"f5", X"03", X"fb", X"03", X"62", X"fa", X"59", X"ff");

begin

process (clk)
  begin
    if rising_edge(clk) then
      dout <= ROM(TO_INTEGER(addr));
    end if;
  end process;

end rtl;
